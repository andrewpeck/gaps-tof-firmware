-- TODO: Need for pulse extension
--         -- make it programmable
-- TODO: Need for alignment
--          -- add inferred SRL16s (prior to the deserializer)
-- TODO: Connect idelays to wishboen
-- TODO: need tx logic
-- TODO: add prbs tx/rx
-- TODO: channel masking
-- TODO: async oversampling? multi-phase clock w/ cd?
--         need to decide if LTMT link carries a clock

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.constants.all;
use work.components.all;
use work.registers.all;
use work.mt_types.all;
use work.ipbus_pkg.all;
use work.types_pkg.all;

entity gaps_mt is
  port(
    --
    clk_i : in std_logic;

    --
    -- eth_rx_d   : in  std_logic_vector (3 downto 0);
    -- eth_rx_dv  : in  std_logic;
    -- eth_rx_clk : in  std_logic;
    -- eth_tx_d   : out std_logic_vector (3 downto 0);
    -- eth_tx_dv  : out std_logic;
    -- eth_tx_clk : out std_logic;

    lt_data_i : in std_logic_vector (NUM_LT_INPUTS-1 downto 0);
    rb_data_o : out std_logic_vector (NUM_RB_OUTPUTS-1 downto 0);
    sump_o : out std_logic
    );
end gaps_mt;

architecture structural of gaps_mt is

  signal locked : std_logic;

  signal clk100, clk200 : std_logic;
  signal clock : std_logic;

  signal event_cnt     : std_logic_vector (EVENTCNTB-1 downto 0);
  signal rst_event_cnt : std_logic := '0';

  -- data/clk delays in units of 78 ps (0-31)
  --  use to align clock/data from a single LT
  signal fine_delays : lt_fine_delays_array_t
    := (others => (others => (others => '0')));
  signal coarse_delays : lt_coarse_delays_array_t
    := (others => (others => (others => '0')));
  signal pulse_stretch : std_logic_vector (3 downto 0)
    := (others => '0');

  signal hits           : channel_array_t;
  signal global_trigger : std_logic;
  signal triggers       : channel_array_t;

  --IPbus
  signal ipb_reset : std_logic;
  signal ipb_clk   : std_logic;
  signal ipb_miso_arr
    : ipb_rbus_array(IPB_SLAVES - 1 downto 0)
    := (others =>
        (ipb_rdata => (others => '0'),
         ipb_ack   => '0',
         ipb_err   => '0'));

  signal ipb_mosi_arr : ipb_wbus_array(IPB_SLAVES - 1 downto 0);

  ------ Register signals begin (this section is generated by generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_MT_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_write_arr       : t_std32_array(REG_MT_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_addresses       : t_std32_array(REG_MT_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_defaults        : t_std32_array(REG_MT_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_MT_NUM_REGS - 1 downto 0) := (others => '0');
    signal regs_write_pulse_arr : std_logic_vector(REG_MT_NUM_REGS - 1 downto 0) := (others => '0');
    signal regs_read_ready_arr  : std_logic_vector(REG_MT_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_MT_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_MT_NUM_REGS - 1 downto 0) := (others => '0');
    -- Connect counter signal declarations
  ------ Register signals end ----------------------------------------------

begin

  clock <= clk100;

  -- take in a global clock, generate system clocks at the correct frequency
  clocking : entity work.clocking
    port map (
      clock_i => clk_i,
      clk100  => clk100,                -- system clock
      clk200  => clk200,                -- 200mhz for iodelay
      locked  => locked                 -- mmcm locked
      );

  -- deserialize and align the inputs
  input_rx : entity work.input_rx
    port map (
      -- system clock
      clk      => clk100, -- logic clock
      clk200   => clk200, -- for idelay

      -- clock and data from lt boards
      clocks_i => (others => clk100),
      data_i   => lt_data_i,

      -- -- idelay settings (in units of 80ps)
      -- clk_delays_i => clk_delays,

      -- sr delay settings (in units of 1 clock cycle)
      fine_delays_i   => fine_delays,
      coarse_delays_i => coarse_delays,

      -- parameter to optionally stretch pulses
      pulse_stretch_i => pulse_stretch,

      -- hit outputs
      hits_o => hits
      );

  -- core trigger logic:
  --   take in a list of hits on channels
  --   return a global OR of the trigger list
  --   and a list of channels to be read out
  trigger : entity work.trigger
    port map (
      -- system clock
      clk => clk100,

      -- hits from input stage (20x16 array of hits)
      hits_i => hits,

      single_hit_en_i => '1', 

      -- ouptut from trigger logic
      global_trigger_o => global_trigger,  -- OR of the trigger menu
      rb_triggers_o    => open,            -- 40 trigger outputs  (1 per rb) 
      triggers_o       => triggers         -- trigger output (320 trigger outputs) 
      );

  -- event counter:
  event_counter : entity work.event_counter
    port map (
      clk              => clock,
      rst_i            => not locked or rst_event_cnt,
      global_trigger_i => global_trigger,
    --trigger_i        => triggers,
      event_count_o    => event_cnt
      );

  sump_o <= global_trigger xor reduce_or(event_cnt);

  -- trg_tx_1: entity work.trg_tx
  --   generic map (
  --     EN_MASK   => EN_MASK,
  --     EVENTCNTB => EVENTCNTB,
  --     MASKCNTB  => MASKCNTB)
  --   port map (
  --     clock       => clock,
  --     reset       => reset,
  --     serial_o    => serial_o,
  --     trg_i       => trg_i,
  --     resync_i    => resync_i,
  --     event_cnt_i => event_cnt_i,
  --     ch_mask_i   => ch_mask_i);

  -- serialize output to the readout boards
  --
  -- output_tx : entity work.output_tx
  --   port map (
  --     clk           => clk,
  --     rst           => not locked,
  --     event_count_i => event_cnt,
  --     trigger_i     => triggers,
  --     trigger_o     => rb_data_o
  --     );

  --===============================================================================================
  --
  --
  -- beyond this is generated by tools/generate_registers.py -- do not edit
  --
  --
  --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave_tmr
        generic map(
           g_ENABLE_TMR           => EN_TMR_IPB_SLAVE_MT,
           g_NUM_REGS             => REG_MT_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_MT_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_MT_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset,
           ipb_clk_i              => ipb_clk,
           ipb_mosi_i             => ipb_mosi_arr(0),
           ipb_miso_o             => ipb_miso_arr(0),
           usr_clk_i              => clock,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"10";
    regs_addresses(1)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"11";
    regs_addresses(2)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"12";
    regs_addresses(3)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"13";
    regs_addresses(4)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"14";
    regs_addresses(5)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"15";
    regs_addresses(6)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"16";
    regs_addresses(7)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"17";
    regs_addresses(8)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"18";
    regs_addresses(9)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"19";
    regs_addresses(10)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"1a";
    regs_addresses(11)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"1b";
    regs_addresses(12)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"1c";
    regs_addresses(13)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"1d";
    regs_addresses(14)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"1e";
    regs_addresses(15)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"1f";
    regs_addresses(16)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"20";
    regs_addresses(17)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"21";
    regs_addresses(18)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"22";
    regs_addresses(19)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"23";
    regs_addresses(20)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"60";
    regs_addresses(21)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"61";
    regs_addresses(22)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"62";
    regs_addresses(23)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"63";
    regs_addresses(24)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"64";
    regs_addresses(25)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"65";
    regs_addresses(26)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"66";
    regs_addresses(27)(REG_MT_ADDRESS_MSB downto REG_MT_ADDRESS_LSB) <= '0' & x"67";

    -- Connect read signals
    regs_read_arr(0)(REG_MT_HIT_COUNTERS_RB0_MSB downto REG_MT_HIT_COUNTERS_RB0_LSB) <= hit_count(0);
    regs_read_arr(1)(REG_MT_HIT_COUNTERS_RB1_MSB downto REG_MT_HIT_COUNTERS_RB1_LSB) <= hit_count(1);
    regs_read_arr(2)(REG_MT_HIT_COUNTERS_RB2_MSB downto REG_MT_HIT_COUNTERS_RB2_LSB) <= hit_count(2);
    regs_read_arr(3)(REG_MT_HIT_COUNTERS_RB3_MSB downto REG_MT_HIT_COUNTERS_RB3_LSB) <= hit_count(3);
    regs_read_arr(4)(REG_MT_HIT_COUNTERS_RB4_MSB downto REG_MT_HIT_COUNTERS_RB4_LSB) <= hit_count(4);
    regs_read_arr(5)(REG_MT_HIT_COUNTERS_RB5_MSB downto REG_MT_HIT_COUNTERS_RB5_LSB) <= hit_count(5);
    regs_read_arr(6)(REG_MT_HIT_COUNTERS_RB6_MSB downto REG_MT_HIT_COUNTERS_RB6_LSB) <= hit_count(6);
    regs_read_arr(7)(REG_MT_HIT_COUNTERS_RB7_MSB downto REG_MT_HIT_COUNTERS_RB7_LSB) <= hit_count(7);
    regs_read_arr(8)(REG_MT_HIT_COUNTERS_RB8_MSB downto REG_MT_HIT_COUNTERS_RB8_LSB) <= hit_count(8);
    regs_read_arr(9)(REG_MT_HIT_COUNTERS_RB9_MSB downto REG_MT_HIT_COUNTERS_RB9_LSB) <= hit_count(9);
    regs_read_arr(10)(REG_MT_HIT_COUNTERS_RB10_MSB downto REG_MT_HIT_COUNTERS_RB10_LSB) <= hit_count(10);
    regs_read_arr(11)(REG_MT_HIT_COUNTERS_RB11_MSB downto REG_MT_HIT_COUNTERS_RB11_LSB) <= hit_count(11);
    regs_read_arr(12)(REG_MT_HIT_COUNTERS_RB12_MSB downto REG_MT_HIT_COUNTERS_RB12_LSB) <= hit_count(12);
    regs_read_arr(13)(REG_MT_HIT_COUNTERS_RB13_MSB downto REG_MT_HIT_COUNTERS_RB13_LSB) <= hit_count(13);
    regs_read_arr(14)(REG_MT_HIT_COUNTERS_RB14_MSB downto REG_MT_HIT_COUNTERS_RB14_LSB) <= hit_count(14);
    regs_read_arr(15)(REG_MT_HIT_COUNTERS_RB15_MSB downto REG_MT_HIT_COUNTERS_RB15_LSB) <= hit_count(15);
    regs_read_arr(16)(REG_MT_HIT_COUNTERS_RB16_MSB downto REG_MT_HIT_COUNTERS_RB16_LSB) <= hit_count(16);
    regs_read_arr(17)(REG_MT_HIT_COUNTERS_RB17_MSB downto REG_MT_HIT_COUNTERS_RB17_LSB) <= hit_count(17);
    regs_read_arr(18)(REG_MT_HIT_COUNTERS_RB18_MSB downto REG_MT_HIT_COUNTERS_RB18_LSB) <= hit_count(18);
    regs_read_arr(19)(REG_MT_HIT_COUNTERS_RB19_MSB downto REG_MT_HIT_COUNTERS_RB19_LSB) <= hit_count(19);
    regs_read_arr(20)(REG_MT_HOG_GLOBAL_DATE_MSB downto REG_MT_HOG_GLOBAL_DATE_LSB) <= GLOBAL_DATE;
    regs_read_arr(21)(REG_MT_HOG_GLOBAL_TIME_MSB downto REG_MT_HOG_GLOBAL_TIME_LSB) <= GLOBAL_TIME;
    regs_read_arr(22)(REG_MT_HOG_GLOBAL_VER_MSB downto REG_MT_HOG_GLOBAL_VER_LSB) <= GLOBAL_VER;
    regs_read_arr(23)(REG_MT_HOG_GLOBAL_SHA_MSB downto REG_MT_HOG_GLOBAL_SHA_LSB) <= GLOBAL_SHA;
    regs_read_arr(24)(REG_MT_HOG_TOP_SHA_MSB downto REG_MT_HOG_TOP_SHA_LSB) <= TOP_SHA;
    regs_read_arr(25)(REG_MT_HOG_TOP_VER_MSB downto REG_MT_HOG_TOP_VER_LSB) <= TOP_VER;
    regs_read_arr(26)(REG_MT_HOG_HOG_SHA_MSB downto REG_MT_HOG_HOG_SHA_LSB) <= HOG_SHA;
    regs_read_arr(27)(REG_MT_HOG_HOG_VER_MSB downto REG_MT_HOG_HOG_VER_LSB) <= HOG_VER;

    -- Connect write signals

    -- Connect write pulse signals

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect counter instances

    COUNTER_MT_HIT_COUNTERS_RB0 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(0)),
        snap_i    => '1',
        count_o   => hit_count(0)
    );


    COUNTER_MT_HIT_COUNTERS_RB1 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(1)),
        snap_i    => '1',
        count_o   => hit_count(1)
    );


    COUNTER_MT_HIT_COUNTERS_RB2 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(2)),
        snap_i    => '1',
        count_o   => hit_count(2)
    );


    COUNTER_MT_HIT_COUNTERS_RB3 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(3)),
        snap_i    => '1',
        count_o   => hit_count(3)
    );


    COUNTER_MT_HIT_COUNTERS_RB4 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(4)),
        snap_i    => '1',
        count_o   => hit_count(4)
    );


    COUNTER_MT_HIT_COUNTERS_RB5 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(5)),
        snap_i    => '1',
        count_o   => hit_count(5)
    );


    COUNTER_MT_HIT_COUNTERS_RB6 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(6)),
        snap_i    => '1',
        count_o   => hit_count(6)
    );


    COUNTER_MT_HIT_COUNTERS_RB7 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(7)),
        snap_i    => '1',
        count_o   => hit_count(7)
    );


    COUNTER_MT_HIT_COUNTERS_RB8 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(8)),
        snap_i    => '1',
        count_o   => hit_count(8)
    );


    COUNTER_MT_HIT_COUNTERS_RB9 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(9)),
        snap_i    => '1',
        count_o   => hit_count(9)
    );


    COUNTER_MT_HIT_COUNTERS_RB10 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(10)),
        snap_i    => '1',
        count_o   => hit_count(10)
    );


    COUNTER_MT_HIT_COUNTERS_RB11 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(11)),
        snap_i    => '1',
        count_o   => hit_count(11)
    );


    COUNTER_MT_HIT_COUNTERS_RB12 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(12)),
        snap_i    => '1',
        count_o   => hit_count(12)
    );


    COUNTER_MT_HIT_COUNTERS_RB13 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(13)),
        snap_i    => '1',
        count_o   => hit_count(13)
    );


    COUNTER_MT_HIT_COUNTERS_RB14 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(14)),
        snap_i    => '1',
        count_o   => hit_count(14)
    );


    COUNTER_MT_HIT_COUNTERS_RB15 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(15)),
        snap_i    => '1',
        count_o   => hit_count(15)
    );


    COUNTER_MT_HIT_COUNTERS_RB16 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(16)),
        snap_i    => '1',
        count_o   => hit_count(16)
    );


    COUNTER_MT_HIT_COUNTERS_RB17 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(17)),
        snap_i    => '1',
        count_o   => hit_count(17)
    );


    COUNTER_MT_HIT_COUNTERS_RB18 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(18)),
        snap_i    => '1',
        count_o   => hit_count(18)
    );


    COUNTER_MT_HIT_COUNTERS_RB19 : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 16
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset,
        en_i      => reduce_or(hits(19)),
        snap_i    => '1',
        count_o   => hit_count(19)
    );


    -- Connect rate instances

    -- Connect read ready signals

    -- Defaults

    -- Define writable regs

--==== Registers end ============================================================================
end structural;
