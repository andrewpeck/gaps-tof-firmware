library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.types_pkg.all;
use work.mt_types.all;
use work.constants.all;
use work.components.all;

entity rb_map is
  port(
    clock         : in  std_logic;
    hit_bitmap_i        : in  channel_bitmask_t := (others => '0');
    rb_ch_bitmap_o : out std_logic_vector (NUM_RBS*8-1 downto 0)
    );
end rb_map;

architecture behavioral of rb_map is
begin

  rb_ch_bitmap_o(0)   <= hit_bitmap_i(0);
  rb_ch_bitmap_o(1)   <= hit_bitmap_i(0);
  rb_ch_bitmap_o(2)   <= hit_bitmap_i(1);
  rb_ch_bitmap_o(3)   <= hit_bitmap_i(1);
  rb_ch_bitmap_o(4)   <= hit_bitmap_i(2);
  rb_ch_bitmap_o(5)   <= hit_bitmap_i(2);
  rb_ch_bitmap_o(6)   <= hit_bitmap_i(3);
  rb_ch_bitmap_o(7)   <= hit_bitmap_i(3);
  rb_ch_bitmap_o(8)   <= hit_bitmap_i(4);
  rb_ch_bitmap_o(9)   <= hit_bitmap_i(4);
  rb_ch_bitmap_o(10)  <= hit_bitmap_i(5);
  rb_ch_bitmap_o(11)  <= hit_bitmap_i(5);
  rb_ch_bitmap_o(12)  <= hit_bitmap_i(6);
  rb_ch_bitmap_o(13)  <= hit_bitmap_i(6);
  rb_ch_bitmap_o(14)  <= hit_bitmap_i(7);
  rb_ch_bitmap_o(15)  <= hit_bitmap_i(7);
  rb_ch_bitmap_o(16)  <= hit_bitmap_i(8);
  rb_ch_bitmap_o(17)  <= hit_bitmap_i(8);
  rb_ch_bitmap_o(18)  <= hit_bitmap_i(9);
  rb_ch_bitmap_o(19)  <= hit_bitmap_i(9);
  rb_ch_bitmap_o(20)  <= hit_bitmap_i(10);
  rb_ch_bitmap_o(21)  <= hit_bitmap_i(10);
  rb_ch_bitmap_o(22)  <= hit_bitmap_i(11);
  rb_ch_bitmap_o(23)  <= hit_bitmap_i(11);
  rb_ch_bitmap_o(24)  <= hit_bitmap_i(12);
  rb_ch_bitmap_o(25)  <= hit_bitmap_i(12);
  rb_ch_bitmap_o(26)  <= hit_bitmap_i(13);
  rb_ch_bitmap_o(27)  <= hit_bitmap_i(13);
  rb_ch_bitmap_o(28)  <= hit_bitmap_i(14);
  rb_ch_bitmap_o(29)  <= hit_bitmap_i(14);
  rb_ch_bitmap_o(30)  <= hit_bitmap_i(15);
  rb_ch_bitmap_o(31)  <= hit_bitmap_i(15);
  rb_ch_bitmap_o(32)  <= hit_bitmap_i(16);
  rb_ch_bitmap_o(33)  <= hit_bitmap_i(16);
  rb_ch_bitmap_o(34)  <= hit_bitmap_i(17);
  rb_ch_bitmap_o(35)  <= hit_bitmap_i(17);
  rb_ch_bitmap_o(36)  <= hit_bitmap_i(18);
  rb_ch_bitmap_o(37)  <= hit_bitmap_i(18);
  rb_ch_bitmap_o(38)  <= hit_bitmap_i(19);
  rb_ch_bitmap_o(39)  <= hit_bitmap_i(19);
  rb_ch_bitmap_o(40)  <= hit_bitmap_i(20);
  rb_ch_bitmap_o(41)  <= hit_bitmap_i(20);
  rb_ch_bitmap_o(42)  <= hit_bitmap_i(21);
  rb_ch_bitmap_o(43)  <= hit_bitmap_i(21);
  rb_ch_bitmap_o(44)  <= hit_bitmap_i(22);
  rb_ch_bitmap_o(45)  <= hit_bitmap_i(22);
  rb_ch_bitmap_o(46)  <= hit_bitmap_i(23);
  rb_ch_bitmap_o(47)  <= hit_bitmap_i(23);
  rb_ch_bitmap_o(48)  <= hit_bitmap_i(24);
  rb_ch_bitmap_o(49)  <= hit_bitmap_i(24);
  rb_ch_bitmap_o(50)  <= hit_bitmap_i(25);
  rb_ch_bitmap_o(51)  <= hit_bitmap_i(25);
  rb_ch_bitmap_o(52)  <= hit_bitmap_i(26);
  rb_ch_bitmap_o(53)  <= hit_bitmap_i(26);
  rb_ch_bitmap_o(54)  <= hit_bitmap_i(27);
  rb_ch_bitmap_o(55)  <= hit_bitmap_i(27);
  rb_ch_bitmap_o(56)  <= hit_bitmap_i(28);
  rb_ch_bitmap_o(57)  <= hit_bitmap_i(28);
  rb_ch_bitmap_o(58)  <= hit_bitmap_i(29);
  rb_ch_bitmap_o(59)  <= hit_bitmap_i(29);
  rb_ch_bitmap_o(60)  <= hit_bitmap_i(30);
  rb_ch_bitmap_o(61)  <= hit_bitmap_i(30);
  rb_ch_bitmap_o(62)  <= hit_bitmap_i(31);
  rb_ch_bitmap_o(63)  <= hit_bitmap_i(31);
  rb_ch_bitmap_o(64)  <= hit_bitmap_i(32);
  rb_ch_bitmap_o(65)  <= hit_bitmap_i(32);
  rb_ch_bitmap_o(66)  <= hit_bitmap_i(33);
  rb_ch_bitmap_o(67)  <= hit_bitmap_i(33);
  rb_ch_bitmap_o(68)  <= hit_bitmap_i(34);
  rb_ch_bitmap_o(69)  <= hit_bitmap_i(34);
  rb_ch_bitmap_o(70)  <= hit_bitmap_i(35);
  rb_ch_bitmap_o(71)  <= hit_bitmap_i(35);
  rb_ch_bitmap_o(72)  <= hit_bitmap_i(36);
  rb_ch_bitmap_o(73)  <= hit_bitmap_i(36);
  rb_ch_bitmap_o(74)  <= hit_bitmap_i(37);
  rb_ch_bitmap_o(75)  <= hit_bitmap_i(37);
  rb_ch_bitmap_o(76)  <= hit_bitmap_i(38);
  rb_ch_bitmap_o(77)  <= hit_bitmap_i(38);
  rb_ch_bitmap_o(78)  <= hit_bitmap_i(39);
  rb_ch_bitmap_o(79)  <= hit_bitmap_i(39);
  rb_ch_bitmap_o(80)  <= hit_bitmap_i(40);
  rb_ch_bitmap_o(81)  <= hit_bitmap_i(40);
  rb_ch_bitmap_o(82)  <= hit_bitmap_i(41);
  rb_ch_bitmap_o(83)  <= hit_bitmap_i(41);
  rb_ch_bitmap_o(84)  <= hit_bitmap_i(42);
  rb_ch_bitmap_o(85)  <= hit_bitmap_i(42);
  rb_ch_bitmap_o(86)  <= hit_bitmap_i(43);
  rb_ch_bitmap_o(87)  <= hit_bitmap_i(43);
  rb_ch_bitmap_o(88)  <= hit_bitmap_i(44);
  rb_ch_bitmap_o(89)  <= hit_bitmap_i(44);
  rb_ch_bitmap_o(90)  <= hit_bitmap_i(45);
  rb_ch_bitmap_o(91)  <= hit_bitmap_i(45);
  rb_ch_bitmap_o(92)  <= hit_bitmap_i(46);
  rb_ch_bitmap_o(93)  <= hit_bitmap_i(46);
  rb_ch_bitmap_o(94)  <= hit_bitmap_i(47);
  rb_ch_bitmap_o(95)  <= hit_bitmap_i(47);
  rb_ch_bitmap_o(96)  <= hit_bitmap_i(48);
  rb_ch_bitmap_o(97)  <= hit_bitmap_i(48);
  rb_ch_bitmap_o(98)  <= hit_bitmap_i(49);
  rb_ch_bitmap_o(99)  <= hit_bitmap_i(49);
  rb_ch_bitmap_o(100) <= hit_bitmap_i(50);
  rb_ch_bitmap_o(101) <= hit_bitmap_i(50);
  rb_ch_bitmap_o(102) <= hit_bitmap_i(51);
  rb_ch_bitmap_o(103) <= hit_bitmap_i(51);
  rb_ch_bitmap_o(104) <= hit_bitmap_i(52);
  rb_ch_bitmap_o(105) <= hit_bitmap_i(52);
  rb_ch_bitmap_o(106) <= hit_bitmap_i(53);
  rb_ch_bitmap_o(107) <= hit_bitmap_i(53);
  rb_ch_bitmap_o(108) <= hit_bitmap_i(54);
  rb_ch_bitmap_o(109) <= hit_bitmap_i(54);
  rb_ch_bitmap_o(110) <= hit_bitmap_i(55);
  rb_ch_bitmap_o(111) <= hit_bitmap_i(55);
  rb_ch_bitmap_o(112) <= hit_bitmap_i(56);
  rb_ch_bitmap_o(113) <= hit_bitmap_i(56);
  rb_ch_bitmap_o(114) <= hit_bitmap_i(57);
  rb_ch_bitmap_o(115) <= hit_bitmap_i(57);
  rb_ch_bitmap_o(116) <= hit_bitmap_i(58);
  rb_ch_bitmap_o(117) <= hit_bitmap_i(58);
  rb_ch_bitmap_o(118) <= hit_bitmap_i(59);
  rb_ch_bitmap_o(119) <= hit_bitmap_i(59);
  rb_ch_bitmap_o(120) <= hit_bitmap_i(60);
  rb_ch_bitmap_o(121) <= hit_bitmap_i(60);
  rb_ch_bitmap_o(122) <= hit_bitmap_i(61);
  rb_ch_bitmap_o(123) <= hit_bitmap_i(61);
  rb_ch_bitmap_o(124) <= hit_bitmap_i(62);
  rb_ch_bitmap_o(125) <= hit_bitmap_i(62);
  rb_ch_bitmap_o(126) <= hit_bitmap_i(63);
  rb_ch_bitmap_o(127) <= hit_bitmap_i(63);
  rb_ch_bitmap_o(128) <= hit_bitmap_i(64);
  rb_ch_bitmap_o(129) <= hit_bitmap_i(64);
  rb_ch_bitmap_o(130) <= hit_bitmap_i(65);
  rb_ch_bitmap_o(131) <= hit_bitmap_i(65);
  rb_ch_bitmap_o(132) <= hit_bitmap_i(66);
  rb_ch_bitmap_o(133) <= hit_bitmap_i(66);
  rb_ch_bitmap_o(134) <= hit_bitmap_i(67);
  rb_ch_bitmap_o(135) <= hit_bitmap_i(67);
  rb_ch_bitmap_o(136) <= hit_bitmap_i(68);
  rb_ch_bitmap_o(137) <= hit_bitmap_i(68);
  rb_ch_bitmap_o(138) <= hit_bitmap_i(69);
  rb_ch_bitmap_o(139) <= hit_bitmap_i(69);
  rb_ch_bitmap_o(140) <= hit_bitmap_i(70);
  rb_ch_bitmap_o(141) <= hit_bitmap_i(70);
  rb_ch_bitmap_o(142) <= hit_bitmap_i(71);
  rb_ch_bitmap_o(143) <= hit_bitmap_i(71);
  rb_ch_bitmap_o(144) <= hit_bitmap_i(72);
  rb_ch_bitmap_o(145) <= hit_bitmap_i(72);
  rb_ch_bitmap_o(146) <= hit_bitmap_i(73);
  rb_ch_bitmap_o(147) <= hit_bitmap_i(73);
  rb_ch_bitmap_o(148) <= hit_bitmap_i(74);
  rb_ch_bitmap_o(149) <= hit_bitmap_i(74);
  rb_ch_bitmap_o(150) <= hit_bitmap_i(75);
  rb_ch_bitmap_o(151) <= hit_bitmap_i(75);
  rb_ch_bitmap_o(152) <= hit_bitmap_i(76);
  rb_ch_bitmap_o(153) <= hit_bitmap_i(76);
  rb_ch_bitmap_o(154) <= hit_bitmap_i(77);
  rb_ch_bitmap_o(155) <= hit_bitmap_i(77);
  rb_ch_bitmap_o(156) <= hit_bitmap_i(78);
  rb_ch_bitmap_o(157) <= hit_bitmap_i(78);
  rb_ch_bitmap_o(158) <= hit_bitmap_i(79);
  rb_ch_bitmap_o(159) <= hit_bitmap_i(79);
  rb_ch_bitmap_o(160) <= hit_bitmap_i(80);
  rb_ch_bitmap_o(161) <= hit_bitmap_i(80);
  rb_ch_bitmap_o(162) <= hit_bitmap_i(81);
  rb_ch_bitmap_o(163) <= hit_bitmap_i(81);
  rb_ch_bitmap_o(164) <= hit_bitmap_i(82);
  rb_ch_bitmap_o(165) <= hit_bitmap_i(82);
  rb_ch_bitmap_o(166) <= hit_bitmap_i(83);
  rb_ch_bitmap_o(167) <= hit_bitmap_i(83);
  rb_ch_bitmap_o(168) <= hit_bitmap_i(84);
  rb_ch_bitmap_o(169) <= hit_bitmap_i(84);
  rb_ch_bitmap_o(170) <= hit_bitmap_i(85);
  rb_ch_bitmap_o(171) <= hit_bitmap_i(85);
  rb_ch_bitmap_o(172) <= hit_bitmap_i(86);
  rb_ch_bitmap_o(173) <= hit_bitmap_i(86);
  rb_ch_bitmap_o(174) <= hit_bitmap_i(87);
  rb_ch_bitmap_o(175) <= hit_bitmap_i(87);
  rb_ch_bitmap_o(176) <= hit_bitmap_i(88);
  rb_ch_bitmap_o(177) <= hit_bitmap_i(88);
  rb_ch_bitmap_o(178) <= hit_bitmap_i(89);
  rb_ch_bitmap_o(179) <= hit_bitmap_i(89);
  rb_ch_bitmap_o(180) <= hit_bitmap_i(90);
  rb_ch_bitmap_o(181) <= hit_bitmap_i(90);
  rb_ch_bitmap_o(182) <= hit_bitmap_i(91);
  rb_ch_bitmap_o(183) <= hit_bitmap_i(91);
  rb_ch_bitmap_o(184) <= hit_bitmap_i(92);
  rb_ch_bitmap_o(185) <= hit_bitmap_i(92);
  rb_ch_bitmap_o(186) <= hit_bitmap_i(93);
  rb_ch_bitmap_o(187) <= hit_bitmap_i(93);
  rb_ch_bitmap_o(188) <= hit_bitmap_i(94);
  rb_ch_bitmap_o(189) <= hit_bitmap_i(94);
  rb_ch_bitmap_o(190) <= hit_bitmap_i(95);
  rb_ch_bitmap_o(191) <= hit_bitmap_i(95);
  rb_ch_bitmap_o(192) <= hit_bitmap_i(96);
  rb_ch_bitmap_o(193) <= hit_bitmap_i(96);
  rb_ch_bitmap_o(194) <= hit_bitmap_i(97);
  rb_ch_bitmap_o(195) <= hit_bitmap_i(97);
  rb_ch_bitmap_o(196) <= hit_bitmap_i(98);
  rb_ch_bitmap_o(197) <= hit_bitmap_i(98);
  rb_ch_bitmap_o(198) <= hit_bitmap_i(99);
  rb_ch_bitmap_o(199) <= hit_bitmap_i(99);
  rb_ch_bitmap_o(200) <= hit_bitmap_i(100);
  rb_ch_bitmap_o(201) <= hit_bitmap_i(100);
  rb_ch_bitmap_o(202) <= hit_bitmap_i(101);
  rb_ch_bitmap_o(203) <= hit_bitmap_i(101);
  rb_ch_bitmap_o(204) <= hit_bitmap_i(102);
  rb_ch_bitmap_o(205) <= hit_bitmap_i(102);
  rb_ch_bitmap_o(206) <= hit_bitmap_i(103);
  rb_ch_bitmap_o(207) <= hit_bitmap_i(103);
  rb_ch_bitmap_o(208) <= hit_bitmap_i(104);
  rb_ch_bitmap_o(209) <= hit_bitmap_i(104);
  rb_ch_bitmap_o(210) <= hit_bitmap_i(105);
  rb_ch_bitmap_o(211) <= hit_bitmap_i(105);
  rb_ch_bitmap_o(212) <= hit_bitmap_i(106);
  rb_ch_bitmap_o(213) <= hit_bitmap_i(106);
  rb_ch_bitmap_o(214) <= hit_bitmap_i(107);
  rb_ch_bitmap_o(215) <= hit_bitmap_i(107);
  rb_ch_bitmap_o(216) <= hit_bitmap_i(108);
  rb_ch_bitmap_o(217) <= hit_bitmap_i(108);
  rb_ch_bitmap_o(218) <= hit_bitmap_i(109);
  rb_ch_bitmap_o(219) <= hit_bitmap_i(109);
  rb_ch_bitmap_o(220) <= hit_bitmap_i(110);
  rb_ch_bitmap_o(221) <= hit_bitmap_i(110);
  rb_ch_bitmap_o(222) <= hit_bitmap_i(111);
  rb_ch_bitmap_o(223) <= hit_bitmap_i(111);
  rb_ch_bitmap_o(224) <= hit_bitmap_i(112);
  rb_ch_bitmap_o(225) <= hit_bitmap_i(112);
  rb_ch_bitmap_o(226) <= hit_bitmap_i(113);
  rb_ch_bitmap_o(227) <= hit_bitmap_i(113);
  rb_ch_bitmap_o(228) <= hit_bitmap_i(114);
  rb_ch_bitmap_o(229) <= hit_bitmap_i(114);
  rb_ch_bitmap_o(230) <= hit_bitmap_i(115);
  rb_ch_bitmap_o(231) <= hit_bitmap_i(115);
  rb_ch_bitmap_o(232) <= hit_bitmap_i(116);
  rb_ch_bitmap_o(233) <= hit_bitmap_i(116);
  rb_ch_bitmap_o(234) <= hit_bitmap_i(117);
  rb_ch_bitmap_o(235) <= hit_bitmap_i(117);
  rb_ch_bitmap_o(236) <= hit_bitmap_i(118);
  rb_ch_bitmap_o(237) <= hit_bitmap_i(118);
  rb_ch_bitmap_o(238) <= hit_bitmap_i(119);
  rb_ch_bitmap_o(239) <= hit_bitmap_i(119);
  rb_ch_bitmap_o(240) <= hit_bitmap_i(120);
  rb_ch_bitmap_o(241) <= hit_bitmap_i(120);
  rb_ch_bitmap_o(242) <= hit_bitmap_i(121);
  rb_ch_bitmap_o(243) <= hit_bitmap_i(121);
  rb_ch_bitmap_o(244) <= hit_bitmap_i(122);
  rb_ch_bitmap_o(245) <= hit_bitmap_i(122);
  rb_ch_bitmap_o(246) <= hit_bitmap_i(123);
  rb_ch_bitmap_o(247) <= hit_bitmap_i(123);
  rb_ch_bitmap_o(248) <= hit_bitmap_i(124);
  rb_ch_bitmap_o(249) <= hit_bitmap_i(124);
  rb_ch_bitmap_o(250) <= hit_bitmap_i(125);
  rb_ch_bitmap_o(251) <= hit_bitmap_i(125);
  rb_ch_bitmap_o(252) <= hit_bitmap_i(126);
  rb_ch_bitmap_o(253) <= hit_bitmap_i(126);
  rb_ch_bitmap_o(254) <= hit_bitmap_i(127);
  rb_ch_bitmap_o(255) <= hit_bitmap_i(127);
  rb_ch_bitmap_o(256) <= hit_bitmap_i(128);
  rb_ch_bitmap_o(257) <= hit_bitmap_i(128);
  rb_ch_bitmap_o(258) <= hit_bitmap_i(129);
  rb_ch_bitmap_o(259) <= hit_bitmap_i(129);
  rb_ch_bitmap_o(260) <= hit_bitmap_i(130);
  rb_ch_bitmap_o(261) <= hit_bitmap_i(130);
  rb_ch_bitmap_o(262) <= hit_bitmap_i(131);
  rb_ch_bitmap_o(263) <= hit_bitmap_i(131);
  rb_ch_bitmap_o(264) <= hit_bitmap_i(132);
  rb_ch_bitmap_o(265) <= hit_bitmap_i(132);
  rb_ch_bitmap_o(266) <= hit_bitmap_i(133);
  rb_ch_bitmap_o(267) <= hit_bitmap_i(133);
  rb_ch_bitmap_o(268) <= hit_bitmap_i(134);
  rb_ch_bitmap_o(269) <= hit_bitmap_i(134);
  rb_ch_bitmap_o(270) <= hit_bitmap_i(135);
  rb_ch_bitmap_o(271) <= hit_bitmap_i(135);
  rb_ch_bitmap_o(272) <= hit_bitmap_i(136);
  rb_ch_bitmap_o(273) <= hit_bitmap_i(136);
  rb_ch_bitmap_o(274) <= hit_bitmap_i(137);
  rb_ch_bitmap_o(275) <= hit_bitmap_i(137);
  rb_ch_bitmap_o(276) <= hit_bitmap_i(138);
  rb_ch_bitmap_o(277) <= hit_bitmap_i(138);
  rb_ch_bitmap_o(278) <= hit_bitmap_i(139);
  rb_ch_bitmap_o(279) <= hit_bitmap_i(139);
  rb_ch_bitmap_o(280) <= hit_bitmap_i(140);
  rb_ch_bitmap_o(281) <= hit_bitmap_i(140);
  rb_ch_bitmap_o(282) <= hit_bitmap_i(141);
  rb_ch_bitmap_o(283) <= hit_bitmap_i(141);
  rb_ch_bitmap_o(284) <= hit_bitmap_i(142);
  rb_ch_bitmap_o(285) <= hit_bitmap_i(142);
  rb_ch_bitmap_o(286) <= hit_bitmap_i(143);
  rb_ch_bitmap_o(287) <= hit_bitmap_i(143);
  rb_ch_bitmap_o(288) <= hit_bitmap_i(144);
  rb_ch_bitmap_o(289) <= hit_bitmap_i(144);
  rb_ch_bitmap_o(290) <= hit_bitmap_i(145);
  rb_ch_bitmap_o(291) <= hit_bitmap_i(145);
  rb_ch_bitmap_o(292) <= hit_bitmap_i(146);
  rb_ch_bitmap_o(293) <= hit_bitmap_i(146);
  rb_ch_bitmap_o(294) <= hit_bitmap_i(147);
  rb_ch_bitmap_o(295) <= hit_bitmap_i(147);
  rb_ch_bitmap_o(296) <= hit_bitmap_i(148);
  rb_ch_bitmap_o(297) <= hit_bitmap_i(148);
  rb_ch_bitmap_o(298) <= hit_bitmap_i(149);
  rb_ch_bitmap_o(299) <= hit_bitmap_i(149);
  rb_ch_bitmap_o(300) <= hit_bitmap_i(150);
  rb_ch_bitmap_o(301) <= hit_bitmap_i(150);
  rb_ch_bitmap_o(302) <= hit_bitmap_i(151);
  rb_ch_bitmap_o(303) <= hit_bitmap_i(151);
  rb_ch_bitmap_o(304) <= hit_bitmap_i(152);
  rb_ch_bitmap_o(305) <= hit_bitmap_i(152);
  rb_ch_bitmap_o(306) <= hit_bitmap_i(153);
  rb_ch_bitmap_o(307) <= hit_bitmap_i(153);
  rb_ch_bitmap_o(308) <= hit_bitmap_i(154);
  rb_ch_bitmap_o(309) <= hit_bitmap_i(154);
  rb_ch_bitmap_o(310) <= hit_bitmap_i(155);
  rb_ch_bitmap_o(311) <= hit_bitmap_i(155);
  rb_ch_bitmap_o(312) <= hit_bitmap_i(156);
  rb_ch_bitmap_o(313) <= hit_bitmap_i(156);
  rb_ch_bitmap_o(314) <= hit_bitmap_i(157);
  rb_ch_bitmap_o(315) <= hit_bitmap_i(157);
  rb_ch_bitmap_o(316) <= hit_bitmap_i(158);
  rb_ch_bitmap_o(317) <= hit_bitmap_i(158);
  rb_ch_bitmap_o(318) <= hit_bitmap_i(159);
  rb_ch_bitmap_o(319) <= hit_bitmap_i(159);
  rb_ch_bitmap_o(320) <= hit_bitmap_i(160);
  rb_ch_bitmap_o(321) <= hit_bitmap_i(160);
  rb_ch_bitmap_o(322) <= hit_bitmap_i(161);
  rb_ch_bitmap_o(323) <= hit_bitmap_i(161);
  rb_ch_bitmap_o(324) <= hit_bitmap_i(162);
  rb_ch_bitmap_o(325) <= hit_bitmap_i(162);
  rb_ch_bitmap_o(326) <= hit_bitmap_i(163);
  rb_ch_bitmap_o(327) <= hit_bitmap_i(163);
  rb_ch_bitmap_o(328) <= hit_bitmap_i(164);
  rb_ch_bitmap_o(329) <= hit_bitmap_i(164);
  rb_ch_bitmap_o(330) <= hit_bitmap_i(165);
  rb_ch_bitmap_o(331) <= hit_bitmap_i(165);
  rb_ch_bitmap_o(332) <= hit_bitmap_i(166);
  rb_ch_bitmap_o(333) <= hit_bitmap_i(166);
  rb_ch_bitmap_o(334) <= hit_bitmap_i(167);
  rb_ch_bitmap_o(335) <= hit_bitmap_i(167);
  rb_ch_bitmap_o(336) <= hit_bitmap_i(168);
  rb_ch_bitmap_o(337) <= hit_bitmap_i(168);
  rb_ch_bitmap_o(338) <= hit_bitmap_i(169);
  rb_ch_bitmap_o(339) <= hit_bitmap_i(169);
  rb_ch_bitmap_o(340) <= hit_bitmap_i(170);
  rb_ch_bitmap_o(341) <= hit_bitmap_i(170);
  rb_ch_bitmap_o(342) <= hit_bitmap_i(171);
  rb_ch_bitmap_o(343) <= hit_bitmap_i(171);
  rb_ch_bitmap_o(344) <= hit_bitmap_i(172);
  rb_ch_bitmap_o(345) <= hit_bitmap_i(172);
  rb_ch_bitmap_o(346) <= hit_bitmap_i(173);
  rb_ch_bitmap_o(347) <= hit_bitmap_i(173);
  rb_ch_bitmap_o(348) <= hit_bitmap_i(174);
  rb_ch_bitmap_o(349) <= hit_bitmap_i(174);
  rb_ch_bitmap_o(350) <= hit_bitmap_i(175);
  rb_ch_bitmap_o(351) <= hit_bitmap_i(175);
  rb_ch_bitmap_o(352) <= hit_bitmap_i(176);
  rb_ch_bitmap_o(353) <= hit_bitmap_i(176);
  rb_ch_bitmap_o(354) <= hit_bitmap_i(177);
  rb_ch_bitmap_o(355) <= hit_bitmap_i(177);
  rb_ch_bitmap_o(356) <= hit_bitmap_i(178);
  rb_ch_bitmap_o(357) <= hit_bitmap_i(178);
  rb_ch_bitmap_o(358) <= hit_bitmap_i(179);
  rb_ch_bitmap_o(359) <= hit_bitmap_i(179);
  rb_ch_bitmap_o(360) <= hit_bitmap_i(180);
  rb_ch_bitmap_o(361) <= hit_bitmap_i(180);
  rb_ch_bitmap_o(362) <= hit_bitmap_i(181);
  rb_ch_bitmap_o(363) <= hit_bitmap_i(181);
  rb_ch_bitmap_o(364) <= hit_bitmap_i(182);
  rb_ch_bitmap_o(365) <= hit_bitmap_i(182);
  rb_ch_bitmap_o(366) <= hit_bitmap_i(183);
  rb_ch_bitmap_o(367) <= hit_bitmap_i(183);
  rb_ch_bitmap_o(368) <= hit_bitmap_i(184);
  rb_ch_bitmap_o(369) <= hit_bitmap_i(184);
  rb_ch_bitmap_o(370) <= hit_bitmap_i(185);
  rb_ch_bitmap_o(371) <= hit_bitmap_i(185);
  rb_ch_bitmap_o(372) <= hit_bitmap_i(186);
  rb_ch_bitmap_o(373) <= hit_bitmap_i(186);
  rb_ch_bitmap_o(374) <= hit_bitmap_i(187);
  rb_ch_bitmap_o(375) <= hit_bitmap_i(187);
  rb_ch_bitmap_o(376) <= hit_bitmap_i(188);
  rb_ch_bitmap_o(377) <= hit_bitmap_i(188);
  rb_ch_bitmap_o(378) <= hit_bitmap_i(189);
  rb_ch_bitmap_o(379) <= hit_bitmap_i(189);
  rb_ch_bitmap_o(380) <= hit_bitmap_i(190);
  rb_ch_bitmap_o(381) <= hit_bitmap_i(190);
  rb_ch_bitmap_o(382) <= hit_bitmap_i(191);
  rb_ch_bitmap_o(383) <= hit_bitmap_i(191);
  rb_ch_bitmap_o(384) <= hit_bitmap_i(192);
  rb_ch_bitmap_o(385) <= hit_bitmap_i(192);
  rb_ch_bitmap_o(386) <= hit_bitmap_i(193);
  rb_ch_bitmap_o(387) <= hit_bitmap_i(193);
  rb_ch_bitmap_o(388) <= hit_bitmap_i(194);
  rb_ch_bitmap_o(389) <= hit_bitmap_i(194);
  rb_ch_bitmap_o(390) <= hit_bitmap_i(195);
  rb_ch_bitmap_o(391) <= hit_bitmap_i(195);
  rb_ch_bitmap_o(392) <= hit_bitmap_i(196);
  rb_ch_bitmap_o(393) <= hit_bitmap_i(196);
  rb_ch_bitmap_o(394) <= hit_bitmap_i(197);
  rb_ch_bitmap_o(395) <= hit_bitmap_i(197);
  rb_ch_bitmap_o(396) <= hit_bitmap_i(198);
  rb_ch_bitmap_o(397) <= hit_bitmap_i(198);
  rb_ch_bitmap_o(398) <= hit_bitmap_i(199);
  rb_ch_bitmap_o(399) <= hit_bitmap_i(199);

end behavioral;
