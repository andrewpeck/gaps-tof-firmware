library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.types_pkg.all;
use work.mt_types.all;
use work.constants.all;
use work.components.all;

entity rb_map is
  port(
    clock          : in  std_logic;
    hits_bitmap_i  : in  channel_bitmask_t := (others => '0');
    rb_ch_bitmap_o : out std_logic_vector (NUM_RBS*8-1 downto 0) := (others => '0') -- 399 downto 0
    );
end rb_map;

architecture behavioral of rb_map is
begin

  -- rb_ch_bitmap_o(399 downto 0) <= hits_bitmap_i(199 downto 0);
  --
  -- this file maps from LTB channels on the right hand side, to readout board
  -- channels on the left hand side.
  --
  -- so e.g. LTB input 0 (DSI1, J1, BIT1) is represented by hits_bitmap_i(0)
  --
  -- the input should be determined by:
  --
  --     CH[0-7] + Harting[0-4]  + DSI[0-5]
  --      * 1         * 8            * 40
  --
  -- the output index should be determined by
  --
  --     CH[0-7]  + Harting Half[0-1] + Harting Number[0-4] + DSI[0-5]
  --      * 1           * 8                  * 16                * 80

  --START: autoinsert mapping

  rb_ch_bitmap_o(  0) <= hits_bitmap_i(  0); -- rb {:board 15, :ch 1} <- ltb {:board 1, :ch 1} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 66, :ltb-num+channel {:board 1, :ch 1}, :rb-num+channel {:board 15, :ch 1}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(  1) <= hits_bitmap_i(  0); -- rb {:board 15, :ch 2} <- ltb {:board 1, :ch 2} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 66, :ltb-num+channel {:board 1, :ch 2}, :rb-num+channel {:board 15, :ch 2}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(  2) <= hits_bitmap_i(  2); -- rb {:board 15, :ch 3} <- ltb {:board 1, :ch 5} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 64, :ltb-num+channel {:board 1, :ch 5}, :rb-num+channel {:board 15, :ch 3}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(  3) <= hits_bitmap_i(  2); -- rb {:board 15, :ch 4} <- ltb {:board 1, :ch 6} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 64, :ltb-num+channel {:board 1, :ch 6}, :rb-num+channel {:board 15, :ch 4}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(  4) <= hits_bitmap_i(  4); -- rb {:board 15, :ch 5} <- ltb {:board 1, :ch 9} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 62, :ltb-num+channel {:board 1, :ch 9}, :rb-num+channel {:board 15, :ch 5}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(  5) <= hits_bitmap_i(  4); -- rb {:board 15, :ch 6} <- ltb {:board 1, :ch 10} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 62, :ltb-num+channel {:board 1, :ch 10}, :rb-num+channel {:board 15, :ch 6}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(  6) <= hits_bitmap_i(  7); -- rb {:board 15, :ch 7} <- ltb {:board 1, :ch 15} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 74, :ltb-num+channel {:board 1, :ch 15}, :rb-num+channel {:board 15, :ch 7}, :dsi-slot 1, :panel-number 8, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(  7) <= hits_bitmap_i(  7); -- rb {:board 15, :ch 8} <- ltb {:board 1, :ch 16} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 74, :ltb-num+channel {:board 1, :ch 16}, :rb-num+channel {:board 15, :ch 8}, :dsi-slot 1, :panel-number 8, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(  8) <= hits_bitmap_i(  1); -- rb {:board 3, :ch 1} <- ltb {:board 1, :ch 3} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 65, :ltb-num+channel {:board 1, :ch 3}, :rb-num+channel {:board 3, :ch 1}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(  9) <= hits_bitmap_i(  1); -- rb {:board 3, :ch 2} <- ltb {:board 1, :ch 4} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 65, :ltb-num+channel {:board 1, :ch 4}, :rb-num+channel {:board 3, :ch 2}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 10) <= hits_bitmap_i(  3); -- rb {:board 3, :ch 3} <- ltb {:board 1, :ch 7} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 63, :ltb-num+channel {:board 1, :ch 7}, :rb-num+channel {:board 3, :ch 3}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 11) <= hits_bitmap_i(  3); -- rb {:board 3, :ch 4} <- ltb {:board 1, :ch 8} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 63, :ltb-num+channel {:board 1, :ch 8}, :rb-num+channel {:board 3, :ch 4}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 12) <= hits_bitmap_i(  5); -- rb {:board 3, :ch 5} <- ltb {:board 1, :ch 11} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 61, :ltb-num+channel {:board 1, :ch 11}, :rb-num+channel {:board 3, :ch 5}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 13) <= hits_bitmap_i(  5); -- rb {:board 3, :ch 6} <- ltb {:board 1, :ch 12} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 61, :ltb-num+channel {:board 1, :ch 12}, :rb-num+channel {:board 3, :ch 6}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 14) <= hits_bitmap_i(  6); -- rb {:board 3, :ch 7} <- ltb {:board 1, :ch 13} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 73, :ltb-num+channel {:board 1, :ch 13}, :rb-num+channel {:board 3, :ch 7}, :dsi-slot 1, :panel-number 8, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 15) <= hits_bitmap_i(  6); -- rb {:board 3, :ch 8} <- ltb {:board 1, :ch 14} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 73, :ltb-num+channel {:board 1, :ch 14}, :rb-num+channel {:board 3, :ch 8}, :dsi-slot 1, :panel-number 8, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 16) <= hits_bitmap_i(  8); -- rb {:board 14, :ch 1} <- ltb {:board 2, :ch 1} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 67, :ltb-num+channel {:board 2, :ch 1}, :rb-num+channel {:board 14, :ch 1}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 17) <= hits_bitmap_i(  8); -- rb {:board 14, :ch 2} <- ltb {:board 2, :ch 2} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 67, :ltb-num+channel {:board 2, :ch 2}, :rb-num+channel {:board 14, :ch 2}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 18) <= hits_bitmap_i( 10); -- rb {:board 14, :ch 3} <- ltb {:board 2, :ch 5} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 69, :ltb-num+channel {:board 2, :ch 5}, :rb-num+channel {:board 14, :ch 3}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 19) <= hits_bitmap_i( 10); -- rb {:board 14, :ch 4} <- ltb {:board 2, :ch 6} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 69, :ltb-num+channel {:board 2, :ch 6}, :rb-num+channel {:board 14, :ch 4}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 20) <= hits_bitmap_i( 12); -- rb {:board 14, :ch 5} <- ltb {:board 2, :ch 9} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 71, :ltb-num+channel {:board 2, :ch 9}, :rb-num+channel {:board 14, :ch 5}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 21) <= hits_bitmap_i( 12); -- rb {:board 14, :ch 6} <- ltb {:board 2, :ch 10} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 71, :ltb-num+channel {:board 2, :ch 10}, :rb-num+channel {:board 14, :ch 6}, :dsi-slot 1, :panel-number 7, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 22) <= hits_bitmap_i( 15); -- rb {:board 14, :ch 7} <- ltb {:board 2, :ch 15} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 92, :ltb-num+channel {:board 2, :ch 15}, :rb-num+channel {:board 14, :ch 7}, :dsi-slot 1, :panel-number 11, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 23) <= hits_bitmap_i( 15); -- rb {:board 14, :ch 8} <- ltb {:board 2, :ch 16} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 92, :ltb-num+channel {:board 2, :ch 16}, :rb-num+channel {:board 14, :ch 8}, :dsi-slot 1, :panel-number 11, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 24) <= hits_bitmap_i(  9); -- rb {:board 32, :ch 1} <- ltb {:board 2, :ch 3} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 68, :ltb-num+channel {:board 2, :ch 3}, :rb-num+channel {:board 32, :ch 1}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 25) <= hits_bitmap_i(  9); -- rb {:board 32, :ch 2} <- ltb {:board 2, :ch 4} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 68, :ltb-num+channel {:board 2, :ch 4}, :rb-num+channel {:board 32, :ch 2}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 26) <= hits_bitmap_i( 11); -- rb {:board 32, :ch 3} <- ltb {:board 2, :ch 7} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 70, :ltb-num+channel {:board 2, :ch 7}, :rb-num+channel {:board 32, :ch 3}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 27) <= hits_bitmap_i( 11); -- rb {:board 32, :ch 4} <- ltb {:board 2, :ch 8} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 70, :ltb-num+channel {:board 2, :ch 8}, :rb-num+channel {:board 32, :ch 4}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 28) <= hits_bitmap_i( 13); -- rb {:board 32, :ch 5} <- ltb {:board 2, :ch 11} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 72, :ltb-num+channel {:board 2, :ch 11}, :rb-num+channel {:board 32, :ch 5}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 29) <= hits_bitmap_i( 13); -- rb {:board 32, :ch 6} <- ltb {:board 2, :ch 12} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 72, :ltb-num+channel {:board 2, :ch 12}, :rb-num+channel {:board 32, :ch 6}, :dsi-slot 1, :panel-number 7, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 30) <= hits_bitmap_i( 14); -- rb {:board 32, :ch 7} <- ltb {:board 2, :ch 13} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 91, :ltb-num+channel {:board 2, :ch 13}, :rb-num+channel {:board 32, :ch 7}, :dsi-slot 1, :panel-number 11, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 31) <= hits_bitmap_i( 14); -- rb {:board 32, :ch 8} <- ltb {:board 2, :ch 14} ::: {:station "umbrella", :ltb-harting 1, :paddle-number 91, :ltb-num+channel {:board 2, :ch 14}, :rb-num+channel {:board 32, :ch 8}, :dsi-slot 1, :panel-number 11, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 32) <= hits_bitmap_i( 16); -- rb {:board 29, :ch 1} <- ltb {:board 3, :ch 1} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 75, :ltb-num+channel {:board 3, :ch 1}, :rb-num+channel {:board 29, :ch 1}, :dsi-slot 1, :panel-number 8, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 33) <= hits_bitmap_i( 16); -- rb {:board 29, :ch 2} <- ltb {:board 3, :ch 2} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 75, :ltb-num+channel {:board 3, :ch 2}, :rb-num+channel {:board 29, :ch 2}, :dsi-slot 1, :panel-number 8, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 34) <= hits_bitmap_i( 18); -- rb {:board 29, :ch 3} <- ltb {:board 3, :ch 5} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 77, :ltb-num+channel {:board 3, :ch 5}, :rb-num+channel {:board 29, :ch 3}, :dsi-slot 1, :panel-number 8, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 35) <= hits_bitmap_i( 18); -- rb {:board 29, :ch 4} <- ltb {:board 3, :ch 6} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 77, :ltb-num+channel {:board 3, :ch 6}, :rb-num+channel {:board 29, :ch 4}, :dsi-slot 1, :panel-number 8, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 36) <= hits_bitmap_i( 21); -- rb {:board 29, :ch 5} <- ltb {:board 3, :ch 11} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 107, :ltb-num+channel {:board 3, :ch 11}, :rb-num+channel {:board 29, :ch 5}, :dsi-slot 1, :panel-number 13, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 37) <= hits_bitmap_i( 21); -- rb {:board 29, :ch 6} <- ltb {:board 3, :ch 12} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 107, :ltb-num+channel {:board 3, :ch 12}, :rb-num+channel {:board 29, :ch 6}, :dsi-slot 1, :panel-number 13, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 38) <= hits_bitmap_i( 23); -- rb {:board 29, :ch 7} <- ltb {:board 3, :ch 15} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 105, :ltb-num+channel {:board 3, :ch 15}, :rb-num+channel {:board 29, :ch 7}, :dsi-slot 1, :panel-number 13, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 39) <= hits_bitmap_i( 23); -- rb {:board 29, :ch 8} <- ltb {:board 3, :ch 16} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 105, :ltb-num+channel {:board 3, :ch 16}, :rb-num+channel {:board 29, :ch 8}, :dsi-slot 1, :panel-number 13, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 40) <= hits_bitmap_i( 17); -- rb {:board 31, :ch 1} <- ltb {:board 3, :ch 3} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 76, :ltb-num+channel {:board 3, :ch 3}, :rb-num+channel {:board 31, :ch 1}, :dsi-slot 1, :panel-number 8, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 41) <= hits_bitmap_i( 17); -- rb {:board 31, :ch 2} <- ltb {:board 3, :ch 4} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 76, :ltb-num+channel {:board 3, :ch 4}, :rb-num+channel {:board 31, :ch 2}, :dsi-slot 1, :panel-number 8, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 42) <= hits_bitmap_i( 19); -- rb {:board 31, :ch 3} <- ltb {:board 3, :ch 7} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 78, :ltb-num+channel {:board 3, :ch 7}, :rb-num+channel {:board 31, :ch 3}, :dsi-slot 1, :panel-number 8, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 43) <= hits_bitmap_i( 19); -- rb {:board 31, :ch 4} <- ltb {:board 3, :ch 8} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 78, :ltb-num+channel {:board 3, :ch 8}, :rb-num+channel {:board 31, :ch 4}, :dsi-slot 1, :panel-number 8, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 44) <= hits_bitmap_i( 20); -- rb {:board 31, :ch 5} <- ltb {:board 3, :ch 9} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 108, :ltb-num+channel {:board 3, :ch 9}, :rb-num+channel {:board 31, :ch 5}, :dsi-slot 1, :panel-number 13, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 45) <= hits_bitmap_i( 20); -- rb {:board 31, :ch 6} <- ltb {:board 3, :ch 10} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 108, :ltb-num+channel {:board 3, :ch 10}, :rb-num+channel {:board 31, :ch 6}, :dsi-slot 1, :panel-number 13, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 46) <= hits_bitmap_i( 22); -- rb {:board 31, :ch 7} <- ltb {:board 3, :ch 13} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 106, :ltb-num+channel {:board 3, :ch 13}, :rb-num+channel {:board 31, :ch 7}, :dsi-slot 1, :panel-number 13, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 47) <= hits_bitmap_i( 22); -- rb {:board 31, :ch 8} <- ltb {:board 3, :ch 14} ::: {:station "umbrella", :ltb-harting 2, :paddle-number 106, :ltb-num+channel {:board 3, :ch 14}, :rb-num+channel {:board 31, :ch 8}, :dsi-slot 1, :panel-number 13, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o( 48) <= hits_bitmap_i( 24); -- rb {:board 13, :ch 1} <- ltb {:board 4, :ch 1} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 93, :ltb-num+channel {:board 4, :ch 1}, :rb-num+channel {:board 13, :ch 1}, :dsi-slot 1, :panel-number 11, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 49) <= hits_bitmap_i( 24); -- rb {:board 13, :ch 2} <- ltb {:board 4, :ch 2} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 93, :ltb-num+channel {:board 4, :ch 2}, :rb-num+channel {:board 13, :ch 2}, :dsi-slot 1, :panel-number 11, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 50) <= hits_bitmap_i( 26); -- rb {:board 13, :ch 3} <- ltb {:board 4, :ch 5} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 95, :ltb-num+channel {:board 4, :ch 5}, :rb-num+channel {:board 13, :ch 3}, :dsi-slot 1, :panel-number 11, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 51) <= hits_bitmap_i( 26); -- rb {:board 13, :ch 4} <- ltb {:board 4, :ch 6} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 95, :ltb-num+channel {:board 4, :ch 6}, :rb-num+channel {:board 13, :ch 4}, :dsi-slot 1, :panel-number 11, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 52) <= hits_bitmap_i( 29); -- rb {:board 13, :ch 5} <- ltb {:board 4, :ch 11} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 89, :ltb-num+channel {:board 4, :ch 11}, :rb-num+channel {:board 13, :ch 5}, :dsi-slot 1, :panel-number 10, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 53) <= hits_bitmap_i( 29); -- rb {:board 13, :ch 6} <- ltb {:board 4, :ch 12} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 89, :ltb-num+channel {:board 4, :ch 12}, :rb-num+channel {:board 13, :ch 6}, :dsi-slot 1, :panel-number 10, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 54) <= hits_bitmap_i( 31); -- rb {:board 13, :ch 7} <- ltb {:board 4, :ch 15} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 87, :ltb-num+channel {:board 4, :ch 15}, :rb-num+channel {:board 13, :ch 7}, :dsi-slot 1, :panel-number 10, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 55) <= hits_bitmap_i( 31); -- rb {:board 13, :ch 8} <- ltb {:board 4, :ch 16} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 87, :ltb-num+channel {:board 4, :ch 16}, :rb-num+channel {:board 13, :ch 8}, :dsi-slot 1, :panel-number 10, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 56) <= hits_bitmap_i( 25); -- rb {:board 35, :ch 1} <- ltb {:board 4, :ch 3} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 94, :ltb-num+channel {:board 4, :ch 3}, :rb-num+channel {:board 35, :ch 1}, :dsi-slot 1, :panel-number 11, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 57) <= hits_bitmap_i( 25); -- rb {:board 35, :ch 2} <- ltb {:board 4, :ch 4} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 94, :ltb-num+channel {:board 4, :ch 4}, :rb-num+channel {:board 35, :ch 2}, :dsi-slot 1, :panel-number 11, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 58) <= hits_bitmap_i( 27); -- rb {:board 35, :ch 3} <- ltb {:board 4, :ch 7} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 96, :ltb-num+channel {:board 4, :ch 7}, :rb-num+channel {:board 35, :ch 3}, :dsi-slot 1, :panel-number 11, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 59) <= hits_bitmap_i( 27); -- rb {:board 35, :ch 4} <- ltb {:board 4, :ch 8} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 96, :ltb-num+channel {:board 4, :ch 8}, :rb-num+channel {:board 35, :ch 4}, :dsi-slot 1, :panel-number 11, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 60) <= hits_bitmap_i( 28); -- rb {:board 35, :ch 5} <- ltb {:board 4, :ch 9} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 90, :ltb-num+channel {:board 4, :ch 9}, :rb-num+channel {:board 35, :ch 5}, :dsi-slot 1, :panel-number 10, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 61) <= hits_bitmap_i( 28); -- rb {:board 35, :ch 6} <- ltb {:board 4, :ch 10} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 90, :ltb-num+channel {:board 4, :ch 10}, :rb-num+channel {:board 35, :ch 6}, :dsi-slot 1, :panel-number 10, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 62) <= hits_bitmap_i( 30); -- rb {:board 35, :ch 7} <- ltb {:board 4, :ch 13} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 88, :ltb-num+channel {:board 4, :ch 13}, :rb-num+channel {:board 35, :ch 7}, :dsi-slot 1, :panel-number 10, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 63) <= hits_bitmap_i( 30); -- rb {:board 35, :ch 8} <- ltb {:board 4, :ch 14} ::: {:station "umbrella", :ltb-harting 3, :paddle-number 88, :ltb-num+channel {:board 4, :ch 14}, :rb-num+channel {:board 35, :ch 8}, :dsi-slot 1, :panel-number 10, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o( 64) <= hits_bitmap_i( 32); -- rb {:board 21, :ch 1} <- ltb {:board 5, :ch 1} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 86, :ltb-num+channel {:board 5, :ch 1}, :rb-num+channel {:board 21, :ch 1}, :dsi-slot 1, :panel-number 10, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 65) <= hits_bitmap_i( 32); -- rb {:board 21, :ch 2} <- ltb {:board 5, :ch 2} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 86, :ltb-num+channel {:board 5, :ch 2}, :rb-num+channel {:board 21, :ch 2}, :dsi-slot 1, :panel-number 10, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 66) <= hits_bitmap_i( 35); -- rb {:board 21, :ch 3} <- ltb {:board 5, :ch 7} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 83, :ltb-num+channel {:board 5, :ch 7}, :rb-num+channel {:board 21, :ch 3}, :dsi-slot 1, :panel-number 9, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 67) <= hits_bitmap_i( 35); -- rb {:board 21, :ch 4} <- ltb {:board 5, :ch 8} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 83, :ltb-num+channel {:board 5, :ch 8}, :rb-num+channel {:board 21, :ch 4}, :dsi-slot 1, :panel-number 9, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 68) <= hits_bitmap_i( 37); -- rb {:board 21, :ch 5} <- ltb {:board 5, :ch 11} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 81, :ltb-num+channel {:board 5, :ch 11}, :rb-num+channel {:board 21, :ch 5}, :dsi-slot 1, :panel-number 9, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 69) <= hits_bitmap_i( 37); -- rb {:board 21, :ch 6} <- ltb {:board 5, :ch 12} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 81, :ltb-num+channel {:board 5, :ch 12}, :rb-num+channel {:board 21, :ch 6}, :dsi-slot 1, :panel-number 9, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 70) <= hits_bitmap_i( 39); -- rb {:board 21, :ch 7} <- ltb {:board 5, :ch 15} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 79, :ltb-num+channel {:board 5, :ch 15}, :rb-num+channel {:board 21, :ch 7}, :dsi-slot 1, :panel-number 9, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 71) <= hits_bitmap_i( 39); -- rb {:board 21, :ch 8} <- ltb {:board 5, :ch 16} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 79, :ltb-num+channel {:board 5, :ch 16}, :rb-num+channel {:board 21, :ch 8}, :dsi-slot 1, :panel-number 9, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 72) <= hits_bitmap_i( 33); -- rb {:board 23, :ch 1} <- ltb {:board 5, :ch 3} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 85, :ltb-num+channel {:board 5, :ch 3}, :rb-num+channel {:board 23, :ch 1}, :dsi-slot 1, :panel-number 10, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 73) <= hits_bitmap_i( 33); -- rb {:board 23, :ch 2} <- ltb {:board 5, :ch 4} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 85, :ltb-num+channel {:board 5, :ch 4}, :rb-num+channel {:board 23, :ch 2}, :dsi-slot 1, :panel-number 10, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 74) <= hits_bitmap_i( 34); -- rb {:board 23, :ch 3} <- ltb {:board 5, :ch 5} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 84, :ltb-num+channel {:board 5, :ch 5}, :rb-num+channel {:board 23, :ch 3}, :dsi-slot 1, :panel-number 9, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 75) <= hits_bitmap_i( 34); -- rb {:board 23, :ch 4} <- ltb {:board 5, :ch 6} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 84, :ltb-num+channel {:board 5, :ch 6}, :rb-num+channel {:board 23, :ch 4}, :dsi-slot 1, :panel-number 9, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 76) <= hits_bitmap_i( 36); -- rb {:board 23, :ch 5} <- ltb {:board 5, :ch 9} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 82, :ltb-num+channel {:board 5, :ch 9}, :rb-num+channel {:board 23, :ch 5}, :dsi-slot 1, :panel-number 9, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 77) <= hits_bitmap_i( 36); -- rb {:board 23, :ch 6} <- ltb {:board 5, :ch 10} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 82, :ltb-num+channel {:board 5, :ch 10}, :rb-num+channel {:board 23, :ch 6}, :dsi-slot 1, :panel-number 9, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 78) <= hits_bitmap_i( 38); -- rb {:board 23, :ch 7} <- ltb {:board 5, :ch 13} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 80, :ltb-num+channel {:board 5, :ch 13}, :rb-num+channel {:board 23, :ch 7}, :dsi-slot 1, :panel-number 9, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 79) <= hits_bitmap_i( 38); -- rb {:board 23, :ch 8} <- ltb {:board 5, :ch 14} ::: {:station "umbrella", :ltb-harting 4, :paddle-number 80, :ltb-num+channel {:board 5, :ch 14}, :rb-num+channel {:board 23, :ch 8}, :dsi-slot 1, :panel-number 9, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o( 80) <= hits_bitmap_i( 40); -- rb {:board 24, :ch 1} <- ltb {:board 6, :ch 1} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 104, :ltb-num+channel {:board 6, :ch 1}, :rb-num+channel {:board 24, :ch 1}, :dsi-slot 2, :panel-number 13, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 81) <= hits_bitmap_i( 40); -- rb {:board 24, :ch 2} <- ltb {:board 6, :ch 2} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 104, :ltb-num+channel {:board 6, :ch 2}, :rb-num+channel {:board 24, :ch 2}, :dsi-slot 2, :panel-number 13, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 82) <= hits_bitmap_i( 43); -- rb {:board 24, :ch 3} <- ltb {:board 6, :ch 7} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 101, :ltb-num+channel {:board 6, :ch 7}, :rb-num+channel {:board 24, :ch 3}, :dsi-slot 2, :panel-number 12, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 83) <= hits_bitmap_i( 43); -- rb {:board 24, :ch 4} <- ltb {:board 6, :ch 8} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 101, :ltb-num+channel {:board 6, :ch 8}, :rb-num+channel {:board 24, :ch 4}, :dsi-slot 2, :panel-number 12, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 84) <= hits_bitmap_i( 45); -- rb {:board 24, :ch 5} <- ltb {:board 6, :ch 11} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 99, :ltb-num+channel {:board 6, :ch 11}, :rb-num+channel {:board 24, :ch 5}, :dsi-slot 2, :panel-number 12, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 85) <= hits_bitmap_i( 45); -- rb {:board 24, :ch 6} <- ltb {:board 6, :ch 12} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 99, :ltb-num+channel {:board 6, :ch 12}, :rb-num+channel {:board 24, :ch 6}, :dsi-slot 2, :panel-number 12, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 86) <= hits_bitmap_i( 47); -- rb {:board 24, :ch 7} <- ltb {:board 6, :ch 15} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 97, :ltb-num+channel {:board 6, :ch 15}, :rb-num+channel {:board 24, :ch 7}, :dsi-slot 2, :panel-number 12, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 87) <= hits_bitmap_i( 47); -- rb {:board 24, :ch 8} <- ltb {:board 6, :ch 16} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 97, :ltb-num+channel {:board 6, :ch 16}, :rb-num+channel {:board 24, :ch 8}, :dsi-slot 2, :panel-number 12, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 88) <= hits_bitmap_i( 41); -- rb {:board 27, :ch 1} <- ltb {:board 6, :ch 3} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 103, :ltb-num+channel {:board 6, :ch 3}, :rb-num+channel {:board 27, :ch 1}, :dsi-slot 2, :panel-number 13, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 89) <= hits_bitmap_i( 41); -- rb {:board 27, :ch 2} <- ltb {:board 6, :ch 4} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 103, :ltb-num+channel {:board 6, :ch 4}, :rb-num+channel {:board 27, :ch 2}, :dsi-slot 2, :panel-number 13, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 90) <= hits_bitmap_i( 42); -- rb {:board 27, :ch 3} <- ltb {:board 6, :ch 5} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 102, :ltb-num+channel {:board 6, :ch 5}, :rb-num+channel {:board 27, :ch 3}, :dsi-slot 2, :panel-number 12, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 91) <= hits_bitmap_i( 42); -- rb {:board 27, :ch 4} <- ltb {:board 6, :ch 6} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 102, :ltb-num+channel {:board 6, :ch 6}, :rb-num+channel {:board 27, :ch 4}, :dsi-slot 2, :panel-number 12, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 92) <= hits_bitmap_i( 44); -- rb {:board 27, :ch 5} <- ltb {:board 6, :ch 9} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 100, :ltb-num+channel {:board 6, :ch 9}, :rb-num+channel {:board 27, :ch 5}, :dsi-slot 2, :panel-number 12, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 93) <= hits_bitmap_i( 44); -- rb {:board 27, :ch 6} <- ltb {:board 6, :ch 10} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 100, :ltb-num+channel {:board 6, :ch 10}, :rb-num+channel {:board 27, :ch 6}, :dsi-slot 2, :panel-number 12, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 94) <= hits_bitmap_i( 46); -- rb {:board 27, :ch 7} <- ltb {:board 6, :ch 13} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 98, :ltb-num+channel {:board 6, :ch 13}, :rb-num+channel {:board 27, :ch 7}, :dsi-slot 2, :panel-number 12, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 95) <= hits_bitmap_i( 46); -- rb {:board 27, :ch 8} <- ltb {:board 6, :ch 14} ::: {:station "umbrella", :ltb-harting 0, :paddle-number 98, :ltb-num+channel {:board 6, :ch 14}, :rb-num+channel {:board 27, :ch 8}, :dsi-slot 2, :panel-number 12, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o( 96) <= hits_bitmap_i( 49); -- rb {:board 40, :ch 1} <- ltb {:board 7, :ch 3} ::: {:station "cortina", :ltb-harting 1, :paddle-number 117, :ltb-num+channel {:board 7, :ch 3}, :rb-num+channel {:board 40, :ch 1}, :dsi-slot 2, :panel-number 14, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o( 97) <= hits_bitmap_i( 49); -- rb {:board 40, :ch 2} <- ltb {:board 7, :ch 4} ::: {:station "cortina", :ltb-harting 1, :paddle-number 117, :ltb-num+channel {:board 7, :ch 4}, :rb-num+channel {:board 40, :ch 2}, :dsi-slot 2, :panel-number 14, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o( 98) <= hits_bitmap_i( 51); -- rb {:board 40, :ch 3} <- ltb {:board 7, :ch 7} ::: {:station "cortina", :ltb-harting 1, :paddle-number 158, :ltb-num+channel {:board 7, :ch 7}, :rb-num+channel {:board 40, :ch 3}, :dsi-slot 2, :panel-number 21, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o( 99) <= hits_bitmap_i( 51); -- rb {:board 40, :ch 4} <- ltb {:board 7, :ch 8} ::: {:station "cortina", :ltb-harting 1, :paddle-number 158, :ltb-num+channel {:board 7, :ch 8}, :rb-num+channel {:board 40, :ch 4}, :dsi-slot 2, :panel-number 21, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(100) <= hits_bitmap_i( 53); -- rb {:board 40, :ch 5} <- ltb {:board 7, :ch 11} ::: {:station "cortina", :ltb-harting 1, :paddle-number 160, :ltb-num+channel {:board 7, :ch 11}, :rb-num+channel {:board 40, :ch 5}, :dsi-slot 2, :panel-number 21, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(101) <= hits_bitmap_i( 53); -- rb {:board 40, :ch 6} <- ltb {:board 7, :ch 12} ::: {:station "cortina", :ltb-harting 1, :paddle-number 160, :ltb-num+channel {:board 7, :ch 12}, :rb-num+channel {:board 40, :ch 6}, :dsi-slot 2, :panel-number 21, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(102) <= hits_bitmap_i( 54); -- rb {:board 40, :ch 7} <- ltb {:board 7, :ch 13} ::: {:station "cube_corner", :ltb-harting 1, :paddle-number 60, :ltb-num+channel {:board 7, :ch 13}, :rb-num+channel {:board 40, :ch 7}, :dsi-slot 2, :panel-number "E-X315", :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(103) <= hits_bitmap_i( 54); -- rb {:board 40, :ch 8} <- ltb {:board 7, :ch 14} ::: {:station "cube_corner", :ltb-harting 1, :paddle-number 60, :ltb-num+channel {:board 7, :ch 14}, :rb-num+channel {:board 40, :ch 8}, :dsi-slot 2, :panel-number "E-X315", :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(104) <= hits_bitmap_i( 48); -- rb {:board 39, :ch 1} <- ltb {:board 7, :ch 1} ::: {:station "cortina", :ltb-harting 1, :paddle-number 116, :ltb-num+channel {:board 7, :ch 1}, :rb-num+channel {:board 39, :ch 1}, :dsi-slot 2, :panel-number 14, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(105) <= hits_bitmap_i( 48); -- rb {:board 39, :ch 2} <- ltb {:board 7, :ch 2} ::: {:station "cortina", :ltb-harting 1, :paddle-number 116, :ltb-num+channel {:board 7, :ch 2}, :rb-num+channel {:board 39, :ch 2}, :dsi-slot 2, :panel-number 14, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(106) <= hits_bitmap_i( 50); -- rb {:board 39, :ch 3} <- ltb {:board 7, :ch 5} ::: {:station "cortina", :ltb-harting 1, :paddle-number 118, :ltb-num+channel {:board 7, :ch 5}, :rb-num+channel {:board 39, :ch 3}, :dsi-slot 2, :panel-number 14, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(107) <= hits_bitmap_i( 50); -- rb {:board 39, :ch 4} <- ltb {:board 7, :ch 6} ::: {:station "cortina", :ltb-harting 1, :paddle-number 118, :ltb-num+channel {:board 7, :ch 6}, :rb-num+channel {:board 39, :ch 4}, :dsi-slot 2, :panel-number 14, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(108) <= hits_bitmap_i( 52); -- rb {:board 39, :ch 5} <- ltb {:board 7, :ch 9} ::: {:station "cortina", :ltb-harting 1, :paddle-number 159, :ltb-num+channel {:board 7, :ch 9}, :rb-num+channel {:board 39, :ch 5}, :dsi-slot 2, :panel-number 21, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(109) <= hits_bitmap_i( 52); -- rb {:board 39, :ch 6} <- ltb {:board 7, :ch 10} ::: {:station "cortina", :ltb-harting 1, :paddle-number 159, :ltb-num+channel {:board 7, :ch 10}, :rb-num+channel {:board 39, :ch 6}, :dsi-slot 2, :panel-number 21, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(110) <= hits_bitmap_i( 55); -- rb {:board 39, :ch 7} <- ltb {:board 7, :ch 15} ::: {:station "cortina", :ltb-harting 1, :paddle-number 148, :ltb-num+channel {:board 7, :ch 15}, :rb-num+channel {:board 39, :ch 7}, :dsi-slot 2, :panel-number 17, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(111) <= hits_bitmap_i( 55); -- rb {:board 39, :ch 8} <- ltb {:board 7, :ch 16} ::: {:station "cortina", :ltb-harting 1, :paddle-number 148, :ltb-num+channel {:board 7, :ch 16}, :rb-num+channel {:board 39, :ch 8}, :dsi-slot 2, :panel-number 17, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o(112) <= hits_bitmap_i( 57); -- rb {:board 25, :ch 1} <- ltb {:board 8, :ch 3} ::: {:station "cube", :ltb-harting 2, :paddle-number 5, :ltb-num+channel {:board 8, :ch 3}, :rb-num+channel {:board 25, :ch 1}, :dsi-slot 2, :panel-number 1, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(113) <= hits_bitmap_i( 57); -- rb {:board 25, :ch 2} <- ltb {:board 8, :ch 4} ::: {:station "cube", :ltb-harting 2, :paddle-number 5, :ltb-num+channel {:board 8, :ch 4}, :rb-num+channel {:board 25, :ch 2}, :dsi-slot 2, :panel-number 1, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(114) <= hits_bitmap_i( 59); -- rb {:board 25, :ch 3} <- ltb {:board 8, :ch 7} ::: {:station "cube", :ltb-harting 2, :paddle-number 3, :ltb-num+channel {:board 8, :ch 7}, :rb-num+channel {:board 25, :ch 3}, :dsi-slot 2, :panel-number 1, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(115) <= hits_bitmap_i( 59); -- rb {:board 25, :ch 4} <- ltb {:board 8, :ch 8} ::: {:station "cube", :ltb-harting 2, :paddle-number 3, :ltb-num+channel {:board 8, :ch 8}, :rb-num+channel {:board 25, :ch 4}, :dsi-slot 2, :panel-number 1, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(116) <= hits_bitmap_i( 61); -- rb {:board 25, :ch 5} <- ltb {:board 8, :ch 11} ::: {:station "cube", :ltb-harting 2, :paddle-number 1, :ltb-num+channel {:board 8, :ch 11}, :rb-num+channel {:board 25, :ch 5}, :dsi-slot 2, :panel-number 1, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(117) <= hits_bitmap_i( 61); -- rb {:board 25, :ch 6} <- ltb {:board 8, :ch 12} ::: {:station "cube", :ltb-harting 2, :paddle-number 1, :ltb-num+channel {:board 8, :ch 12}, :rb-num+channel {:board 25, :ch 6}, :dsi-slot 2, :panel-number 1, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(118) <= hits_bitmap_i( 63); -- rb {:board 25, :ch 7} <- ltb {:board 8, :ch 15} ::: {:station "cube", :ltb-harting 2, :paddle-number 26, :ltb-num+channel {:board 8, :ch 15}, :rb-num+channel {:board 25, :ch 7}, :dsi-slot 2, :panel-number 3, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(119) <= hits_bitmap_i( 63); -- rb {:board 25, :ch 8} <- ltb {:board 8, :ch 16} ::: {:station "cube", :ltb-harting 2, :paddle-number 26, :ltb-num+channel {:board 8, :ch 16}, :rb-num+channel {:board 25, :ch 8}, :dsi-slot 2, :panel-number 3, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(120) <= hits_bitmap_i( 56); -- rb {:board 16, :ch 1} <- ltb {:board 8, :ch 1} ::: {:station "cube", :ltb-harting 2, :paddle-number 6, :ltb-num+channel {:board 8, :ch 1}, :rb-num+channel {:board 16, :ch 1}, :dsi-slot 2, :panel-number 1, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(121) <= hits_bitmap_i( 56); -- rb {:board 16, :ch 2} <- ltb {:board 8, :ch 2} ::: {:station "cube", :ltb-harting 2, :paddle-number 6, :ltb-num+channel {:board 8, :ch 2}, :rb-num+channel {:board 16, :ch 2}, :dsi-slot 2, :panel-number 1, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(122) <= hits_bitmap_i( 58); -- rb {:board 16, :ch 3} <- ltb {:board 8, :ch 5} ::: {:station "cube", :ltb-harting 2, :paddle-number 4, :ltb-num+channel {:board 8, :ch 5}, :rb-num+channel {:board 16, :ch 3}, :dsi-slot 2, :panel-number 1, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(123) <= hits_bitmap_i( 58); -- rb {:board 16, :ch 4} <- ltb {:board 8, :ch 6} ::: {:station "cube", :ltb-harting 2, :paddle-number 4, :ltb-num+channel {:board 8, :ch 6}, :rb-num+channel {:board 16, :ch 4}, :dsi-slot 2, :panel-number 1, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(124) <= hits_bitmap_i( 60); -- rb {:board 16, :ch 5} <- ltb {:board 8, :ch 9} ::: {:station "cube", :ltb-harting 2, :paddle-number 2, :ltb-num+channel {:board 8, :ch 9}, :rb-num+channel {:board 16, :ch 5}, :dsi-slot 2, :panel-number 1, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(125) <= hits_bitmap_i( 60); -- rb {:board 16, :ch 6} <- ltb {:board 8, :ch 10} ::: {:station "cube", :ltb-harting 2, :paddle-number 2, :ltb-num+channel {:board 8, :ch 10}, :rb-num+channel {:board 16, :ch 6}, :dsi-slot 2, :panel-number 1, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(126) <= hits_bitmap_i( 62); -- rb {:board 16, :ch 7} <- ltb {:board 8, :ch 13} ::: {:station "cube", :ltb-harting 2, :paddle-number 25, :ltb-num+channel {:board 8, :ch 13}, :rb-num+channel {:board 16, :ch 7}, :dsi-slot 2, :panel-number 3, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(127) <= hits_bitmap_i( 62); -- rb {:board 16, :ch 8} <- ltb {:board 8, :ch 14} ::: {:station "cube", :ltb-harting 2, :paddle-number 25, :ltb-num+channel {:board 8, :ch 14}, :rb-num+channel {:board 16, :ch 8}, :dsi-slot 2, :panel-number 3, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(128) <= hits_bitmap_i( 64); -- rb {:board 46, :ch 1} <- ltb {:board 9, :ch 1} ::: {:station "cube", :ltb-harting 3, :paddle-number 32, :ltb-num+channel {:board 9, :ch 1}, :rb-num+channel {:board 46, :ch 1}, :dsi-slot 2, :panel-number 3, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(129) <= hits_bitmap_i( 64); -- rb {:board 46, :ch 2} <- ltb {:board 9, :ch 2} ::: {:station "cube", :ltb-harting 3, :paddle-number 32, :ltb-num+channel {:board 9, :ch 2}, :rb-num+channel {:board 46, :ch 2}, :dsi-slot 2, :panel-number 3, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(130) <= hits_bitmap_i( 66); -- rb {:board 46, :ch 3} <- ltb {:board 9, :ch 5} ::: {:station "cube", :ltb-harting 3, :paddle-number 30, :ltb-num+channel {:board 9, :ch 5}, :rb-num+channel {:board 46, :ch 3}, :dsi-slot 2, :panel-number 3, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(131) <= hits_bitmap_i( 66); -- rb {:board 46, :ch 4} <- ltb {:board 9, :ch 6} ::: {:station "cube", :ltb-harting 3, :paddle-number 30, :ltb-num+channel {:board 9, :ch 6}, :rb-num+channel {:board 46, :ch 4}, :dsi-slot 2, :panel-number 3, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(132) <= hits_bitmap_i( 68); -- rb {:board 46, :ch 5} <- ltb {:board 9, :ch 9} ::: {:station "cube", :ltb-harting 3, :paddle-number 28, :ltb-num+channel {:board 9, :ch 9}, :rb-num+channel {:board 46, :ch 5}, :dsi-slot 2, :panel-number 3, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(133) <= hits_bitmap_i( 68); -- rb {:board 46, :ch 6} <- ltb {:board 9, :ch 10} ::: {:station "cube", :ltb-harting 3, :paddle-number 28, :ltb-num+channel {:board 9, :ch 10}, :rb-num+channel {:board 46, :ch 6}, :dsi-slot 2, :panel-number 3, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(134) <= hits_bitmap_i( 70); -- rb {:board 46, :ch 7} <- ltb {:board 9, :ch 13} ::: {:station "cortina", :ltb-harting 3, :paddle-number 110, :ltb-num+channel {:board 9, :ch 13}, :rb-num+channel {:board 46, :ch 7}, :dsi-slot 2, :panel-number 14, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(135) <= hits_bitmap_i( 70); -- rb {:board 46, :ch 8} <- ltb {:board 9, :ch 14} ::: {:station "cortina", :ltb-harting 3, :paddle-number 110, :ltb-num+channel {:board 9, :ch 14}, :rb-num+channel {:board 46, :ch 8}, :dsi-slot 2, :panel-number 14, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(136) <= hits_bitmap_i( 65); -- rb {:board 8, :ch 1} <- ltb {:board 9, :ch 3} ::: {:station "cube", :ltb-harting 3, :paddle-number 31, :ltb-num+channel {:board 9, :ch 3}, :rb-num+channel {:board 8, :ch 1}, :dsi-slot 2, :panel-number 3, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(137) <= hits_bitmap_i( 65); -- rb {:board 8, :ch 2} <- ltb {:board 9, :ch 4} ::: {:station "cube", :ltb-harting 3, :paddle-number 31, :ltb-num+channel {:board 9, :ch 4}, :rb-num+channel {:board 8, :ch 2}, :dsi-slot 2, :panel-number 3, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(138) <= hits_bitmap_i( 67); -- rb {:board 8, :ch 3} <- ltb {:board 9, :ch 7} ::: {:station "cube", :ltb-harting 3, :paddle-number 29, :ltb-num+channel {:board 9, :ch 7}, :rb-num+channel {:board 8, :ch 3}, :dsi-slot 2, :panel-number 3, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(139) <= hits_bitmap_i( 67); -- rb {:board 8, :ch 4} <- ltb {:board 9, :ch 8} ::: {:station "cube", :ltb-harting 3, :paddle-number 29, :ltb-num+channel {:board 9, :ch 8}, :rb-num+channel {:board 8, :ch 4}, :dsi-slot 2, :panel-number 3, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(140) <= hits_bitmap_i( 69); -- rb {:board 8, :ch 5} <- ltb {:board 9, :ch 11} ::: {:station "cube", :ltb-harting 3, :paddle-number 27, :ltb-num+channel {:board 9, :ch 11}, :rb-num+channel {:board 8, :ch 5}, :dsi-slot 2, :panel-number 3, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(141) <= hits_bitmap_i( 69); -- rb {:board 8, :ch 6} <- ltb {:board 9, :ch 12} ::: {:station "cube", :ltb-harting 3, :paddle-number 27, :ltb-num+channel {:board 9, :ch 12}, :rb-num+channel {:board 8, :ch 6}, :dsi-slot 2, :panel-number 3, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(142) <= hits_bitmap_i( 71); -- rb {:board 8, :ch 7} <- ltb {:board 9, :ch 15} ::: {:station "cortina", :ltb-harting 3, :paddle-number 109, :ltb-num+channel {:board 9, :ch 15}, :rb-num+channel {:board 8, :ch 7}, :dsi-slot 2, :panel-number 14, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(143) <= hits_bitmap_i( 71); -- rb {:board 8, :ch 8} <- ltb {:board 9, :ch 16} ::: {:station "cortina", :ltb-harting 3, :paddle-number 109, :ltb-num+channel {:board 9, :ch 16}, :rb-num+channel {:board 8, :ch 8}, :dsi-slot 2, :panel-number 14, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(144) <= hits_bitmap_i( 72); -- rb {:board 11, :ch 1} <- ltb {:board 10, :ch 1} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 13, :ltb-num+channel {:board 10, :ch 1}, :rb-num+channel {:board 11, :ch 1}, :dsi-slot 2, :panel-number 2, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(145) <= hits_bitmap_i( 72); -- rb {:board 11, :ch 2} <- ltb {:board 10, :ch 2} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 13, :ltb-num+channel {:board 10, :ch 2}, :rb-num+channel {:board 11, :ch 2}, :dsi-slot 2, :panel-number 2, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(146) <= hits_bitmap_i( 74); -- rb {:board 11, :ch 3} <- ltb {:board 10, :ch 5} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 15, :ltb-num+channel {:board 10, :ch 5}, :rb-num+channel {:board 11, :ch 3}, :dsi-slot 2, :panel-number 2, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(147) <= hits_bitmap_i( 74); -- rb {:board 11, :ch 4} <- ltb {:board 10, :ch 6} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 15, :ltb-num+channel {:board 10, :ch 6}, :rb-num+channel {:board 11, :ch 4}, :dsi-slot 2, :panel-number 2, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(148) <= hits_bitmap_i( 76); -- rb {:board 11, :ch 5} <- ltb {:board 10, :ch 9} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 17, :ltb-num+channel {:board 10, :ch 9}, :rb-num+channel {:board 11, :ch 5}, :dsi-slot 2, :panel-number 2, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(149) <= hits_bitmap_i( 76); -- rb {:board 11, :ch 6} <- ltb {:board 10, :ch 10} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 17, :ltb-num+channel {:board 10, :ch 10}, :rb-num+channel {:board 11, :ch 6}, :dsi-slot 2, :panel-number 2, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(150) <= hits_bitmap_i( 78); -- rb {:board 11, :ch 7} <- ltb {:board 10, :ch 13} ::: {:station "cortina", :ltb-harting 4, :paddle-number 112, :ltb-num+channel {:board 10, :ch 13}, :rb-num+channel {:board 11, :ch 7}, :dsi-slot 2, :panel-number 14, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(151) <= hits_bitmap_i( 78); -- rb {:board 11, :ch 8} <- ltb {:board 10, :ch 14} ::: {:station "cortina", :ltb-harting 4, :paddle-number 112, :ltb-num+channel {:board 10, :ch 14}, :rb-num+channel {:board 11, :ch 8}, :dsi-slot 2, :panel-number 14, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(152) <= hits_bitmap_i( 73); -- rb {:board 1, :ch 1} <- ltb {:board 10, :ch 3} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 14, :ltb-num+channel {:board 10, :ch 3}, :rb-num+channel {:board 1, :ch 1}, :dsi-slot 2, :panel-number 2, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(153) <= hits_bitmap_i( 73); -- rb {:board 1, :ch 2} <- ltb {:board 10, :ch 4} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 14, :ltb-num+channel {:board 10, :ch 4}, :rb-num+channel {:board 1, :ch 2}, :dsi-slot 2, :panel-number 2, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(154) <= hits_bitmap_i( 75); -- rb {:board 1, :ch 3} <- ltb {:board 10, :ch 7} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 16, :ltb-num+channel {:board 10, :ch 7}, :rb-num+channel {:board 1, :ch 3}, :dsi-slot 2, :panel-number 2, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(155) <= hits_bitmap_i( 75); -- rb {:board 1, :ch 4} <- ltb {:board 10, :ch 8} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 16, :ltb-num+channel {:board 10, :ch 8}, :rb-num+channel {:board 1, :ch 4}, :dsi-slot 2, :panel-number 2, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(156) <= hits_bitmap_i( 77); -- rb {:board 1, :ch 5} <- ltb {:board 10, :ch 11} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 18, :ltb-num+channel {:board 10, :ch 11}, :rb-num+channel {:board 1, :ch 5}, :dsi-slot 2, :panel-number 2, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(157) <= hits_bitmap_i( 77); -- rb {:board 1, :ch 6} <- ltb {:board 10, :ch 12} ::: {:station "cube_bot", :ltb-harting 4, :paddle-number 18, :ltb-num+channel {:board 10, :ch 12}, :rb-num+channel {:board 1, :ch 6}, :dsi-slot 2, :panel-number 2, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(158) <= hits_bitmap_i( 79); -- rb {:board 1, :ch 7} <- ltb {:board 10, :ch 15} ::: {:station "cortina", :ltb-harting 4, :paddle-number 111, :ltb-num+channel {:board 10, :ch 15}, :rb-num+channel {:board 1, :ch 7}, :dsi-slot 2, :panel-number 14, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(159) <= hits_bitmap_i( 79); -- rb {:board 1, :ch 8} <- ltb {:board 10, :ch 16} ::: {:station "cortina", :ltb-harting 4, :paddle-number 111, :ltb-num+channel {:board 10, :ch 16}, :rb-num+channel {:board 1, :ch 8}, :dsi-slot 2, :panel-number 14, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(160) <= hits_bitmap_i( 81); -- rb {:board 42, :ch 1} <- ltb {:board 11, :ch 3} ::: {:station "cube_corner", :ltb-harting 0, :paddle-number 57, :ltb-num+channel {:board 11, :ch 3}, :rb-num+channel {:board 42, :ch 1}, :dsi-slot 3, :panel-number "E-X045", :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(161) <= hits_bitmap_i( 81); -- rb {:board 42, :ch 2} <- ltb {:board 11, :ch 4} ::: {:station "cube_corner", :ltb-harting 0, :paddle-number 57, :ltb-num+channel {:board 11, :ch 4}, :rb-num+channel {:board 42, :ch 2}, :dsi-slot 3, :panel-number "E-X045", :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(162) <= hits_bitmap_i( 85); -- rb {:board 42, :ch 3} <- ltb {:board 11, :ch 11} ::: {:station "cortina", :ltb-harting 0, :paddle-number 149, :ltb-num+channel {:board 11, :ch 11}, :rb-num+channel {:board 42, :ch 3}, :dsi-slot 3, :panel-number 18, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(163) <= hits_bitmap_i( 85); -- rb {:board 42, :ch 4} <- ltb {:board 11, :ch 12} ::: {:station "cortina", :ltb-harting 0, :paddle-number 149, :ltb-num+channel {:board 11, :ch 12}, :rb-num+channel {:board 42, :ch 4}, :dsi-slot 3, :panel-number 18, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(164) <= hits_bitmap_i( 86); -- rb {:board 42, :ch 5} <- ltb {:board 11, :ch 13} ::: {:station "cortina", :ltb-harting 0, :paddle-number 150, :ltb-num+channel {:board 11, :ch 13}, :rb-num+channel {:board 42, :ch 5}, :dsi-slot 3, :panel-number 18, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(165) <= hits_bitmap_i( 86); -- rb {:board 42, :ch 6} <- ltb {:board 11, :ch 14} ::: {:station "cortina", :ltb-harting 0, :paddle-number 150, :ltb-num+channel {:board 11, :ch 14}, :rb-num+channel {:board 42, :ch 6}, :dsi-slot 3, :panel-number 18, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(166) <= hits_bitmap_i( 87); -- rb {:board 42, :ch 7} <- ltb {:board 11, :ch 15} ::: {:station "cortina", :ltb-harting 0, :paddle-number 151, :ltb-num+channel {:board 11, :ch 15}, :rb-num+channel {:board 42, :ch 7}, :dsi-slot 3, :panel-number 18, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(167) <= hits_bitmap_i( 87); -- rb {:board 42, :ch 8} <- ltb {:board 11, :ch 16} ::: {:station "cortina", :ltb-harting 0, :paddle-number 151, :ltb-num+channel {:board 11, :ch 16}, :rb-num+channel {:board 42, :ch 8}, :dsi-slot 3, :panel-number 18, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(168) <= hits_bitmap_i( 80); -- rb {:board 41, :ch 1} <- ltb {:board 11, :ch 1} ::: {:station "cortina", :ltb-harting 0, :paddle-number 128, :ltb-num+channel {:board 11, :ch 1}, :rb-num+channel {:board 41, :ch 1}, :dsi-slot 3, :panel-number 15, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(169) <= hits_bitmap_i( 80); -- rb {:board 41, :ch 2} <- ltb {:board 11, :ch 2} ::: {:station "cortina", :ltb-harting 0, :paddle-number 128, :ltb-num+channel {:board 11, :ch 2}, :rb-num+channel {:board 41, :ch 2}, :dsi-slot 3, :panel-number 15, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(170) <= hits_bitmap_i( 82); -- rb {:board 41, :ch 3} <- ltb {:board 11, :ch 5} ::: {:station "cortina", :ltb-harting 0, :paddle-number 115, :ltb-num+channel {:board 11, :ch 5}, :rb-num+channel {:board 41, :ch 3}, :dsi-slot 3, :panel-number 14, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(171) <= hits_bitmap_i( 82); -- rb {:board 41, :ch 4} <- ltb {:board 11, :ch 6} ::: {:station "cortina", :ltb-harting 0, :paddle-number 115, :ltb-num+channel {:board 11, :ch 6}, :rb-num+channel {:board 41, :ch 4}, :dsi-slot 3, :panel-number 14, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(172) <= hits_bitmap_i( 83); -- rb {:board 41, :ch 5} <- ltb {:board 11, :ch 7} ::: {:station "cortina", :ltb-harting 0, :paddle-number 114, :ltb-num+channel {:board 11, :ch 7}, :rb-num+channel {:board 41, :ch 5}, :dsi-slot 3, :panel-number 14, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(173) <= hits_bitmap_i( 83); -- rb {:board 41, :ch 6} <- ltb {:board 11, :ch 8} ::: {:station "cortina", :ltb-harting 0, :paddle-number 114, :ltb-num+channel {:board 11, :ch 8}, :rb-num+channel {:board 41, :ch 6}, :dsi-slot 3, :panel-number 14, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(174) <= hits_bitmap_i( 84); -- rb {:board 41, :ch 7} <- ltb {:board 11, :ch 9} ::: {:station "cortina", :ltb-harting 0, :paddle-number 113, :ltb-num+channel {:board 11, :ch 9}, :rb-num+channel {:board 41, :ch 7}, :dsi-slot 3, :panel-number 14, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(175) <= hits_bitmap_i( 84); -- rb {:board 41, :ch 8} <- ltb {:board 11, :ch 10} ::: {:station "cortina", :ltb-harting 0, :paddle-number 113, :ltb-num+channel {:board 11, :ch 10}, :rb-num+channel {:board 41, :ch 8}, :dsi-slot 3, :panel-number 14, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(176) <= hits_bitmap_i( 88); -- rb {:board 19, :ch 1} <- ltb {:board 12, :ch 1} ::: {:station "cube", :ltb-harting 1, :paddle-number 40, :ltb-num+channel {:board 12, :ch 1}, :rb-num+channel {:board 19, :ch 1}, :dsi-slot 3, :panel-number 4, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(177) <= hits_bitmap_i( 88); -- rb {:board 19, :ch 2} <- ltb {:board 12, :ch 2} ::: {:station "cube", :ltb-harting 1, :paddle-number 40, :ltb-num+channel {:board 12, :ch 2}, :rb-num+channel {:board 19, :ch 2}, :dsi-slot 3, :panel-number 4, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(178) <= hits_bitmap_i( 89); -- rb {:board 19, :ch 3} <- ltb {:board 12, :ch 3} ::: {:station "cube", :ltb-harting 1, :paddle-number 38, :ltb-num+channel {:board 12, :ch 3}, :rb-num+channel {:board 19, :ch 3}, :dsi-slot 3, :panel-number 4, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(179) <= hits_bitmap_i( 89); -- rb {:board 19, :ch 4} <- ltb {:board 12, :ch 4} ::: {:station "cube", :ltb-harting 1, :paddle-number 38, :ltb-num+channel {:board 12, :ch 4}, :rb-num+channel {:board 19, :ch 4}, :dsi-slot 3, :panel-number 4, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(180) <= hits_bitmap_i( 90); -- rb {:board 19, :ch 5} <- ltb {:board 12, :ch 5} ::: {:station "cube", :ltb-harting 1, :paddle-number 36, :ltb-num+channel {:board 12, :ch 5}, :rb-num+channel {:board 19, :ch 5}, :dsi-slot 3, :panel-number 4, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(181) <= hits_bitmap_i( 90); -- rb {:board 19, :ch 6} <- ltb {:board 12, :ch 6} ::: {:station "cube", :ltb-harting 1, :paddle-number 36, :ltb-num+channel {:board 12, :ch 6}, :rb-num+channel {:board 19, :ch 6}, :dsi-slot 3, :panel-number 4, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(182) <= hits_bitmap_i( 91); -- rb {:board 19, :ch 7} <- ltb {:board 12, :ch 7} ::: {:station "cube", :ltb-harting 1, :paddle-number 34, :ltb-num+channel {:board 12, :ch 7}, :rb-num+channel {:board 19, :ch 7}, :dsi-slot 3, :panel-number 4, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(183) <= hits_bitmap_i( 91); -- rb {:board 19, :ch 8} <- ltb {:board 12, :ch 8} ::: {:station "cube", :ltb-harting 1, :paddle-number 34, :ltb-num+channel {:board 12, :ch 8}, :rb-num+channel {:board 19, :ch 8}, :dsi-slot 3, :panel-number 4, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(184) <= hits_bitmap_i( 95); -- rb {:board 20, :ch 1} <- ltb {:board 12, :ch 15} ::: {:station "cube", :ltb-harting 1, :paddle-number 39, :ltb-num+channel {:board 12, :ch 15}, :rb-num+channel {:board 20, :ch 1}, :dsi-slot 3, :panel-number 4, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(185) <= hits_bitmap_i( 95); -- rb {:board 20, :ch 2} <- ltb {:board 12, :ch 16} ::: {:station "cube", :ltb-harting 1, :paddle-number 39, :ltb-num+channel {:board 12, :ch 16}, :rb-num+channel {:board 20, :ch 2}, :dsi-slot 3, :panel-number 4, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(186) <= hits_bitmap_i( 94); -- rb {:board 20, :ch 3} <- ltb {:board 12, :ch 13} ::: {:station "cube", :ltb-harting 1, :paddle-number 37, :ltb-num+channel {:board 12, :ch 13}, :rb-num+channel {:board 20, :ch 3}, :dsi-slot 3, :panel-number 4, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(187) <= hits_bitmap_i( 94); -- rb {:board 20, :ch 4} <- ltb {:board 12, :ch 14} ::: {:station "cube", :ltb-harting 1, :paddle-number 37, :ltb-num+channel {:board 12, :ch 14}, :rb-num+channel {:board 20, :ch 4}, :dsi-slot 3, :panel-number 4, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(188) <= hits_bitmap_i( 93); -- rb {:board 20, :ch 5} <- ltb {:board 12, :ch 11} ::: {:station "cube", :ltb-harting 1, :paddle-number 35, :ltb-num+channel {:board 12, :ch 11}, :rb-num+channel {:board 20, :ch 5}, :dsi-slot 3, :panel-number 4, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(189) <= hits_bitmap_i( 93); -- rb {:board 20, :ch 6} <- ltb {:board 12, :ch 12} ::: {:station "cube", :ltb-harting 1, :paddle-number 35, :ltb-num+channel {:board 12, :ch 12}, :rb-num+channel {:board 20, :ch 6}, :dsi-slot 3, :panel-number 4, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(190) <= hits_bitmap_i( 92); -- rb {:board 20, :ch 7} <- ltb {:board 12, :ch 9} ::: {:station "cube", :ltb-harting 1, :paddle-number 33, :ltb-num+channel {:board 12, :ch 9}, :rb-num+channel {:board 20, :ch 7}, :dsi-slot 3, :panel-number 4, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(191) <= hits_bitmap_i( 92); -- rb {:board 20, :ch 8} <- ltb {:board 12, :ch 10} ::: {:station "cube", :ltb-harting 1, :paddle-number 33, :ltb-num+channel {:board 12, :ch 10}, :rb-num+channel {:board 20, :ch 8}, :dsi-slot 3, :panel-number 4, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(192) <= hits_bitmap_i( 96); -- rb {:board 18, :ch 1} <- ltb {:board 13, :ch 1} ::: {:station "cortina", :ltb-harting 2, :paddle-number 152, :ltb-num+channel {:board 13, :ch 1}, :rb-num+channel {:board 18, :ch 1}, :dsi-slot 3, :panel-number 19, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(193) <= hits_bitmap_i(101); -- rb {:board 18, :ch 2} <- ltb {:board 13, :ch 12} ::: {:station "cortina", :ltb-harting 2, :paddle-number 152, :ltb-num+channel {:board 13, :ch 12}, :rb-num+channel {:board 18, :ch 2}, :dsi-slot 3, :panel-number 19, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(194) <= hits_bitmap_i( 97); -- rb {:board 18, :ch 3} <- ltb {:board 13, :ch 3} ::: {:station "cortina", :ltb-harting 2, :paddle-number 153, :ltb-num+channel {:board 13, :ch 3}, :rb-num+channel {:board 18, :ch 3}, :dsi-slot 3, :panel-number 19, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(195) <= hits_bitmap_i( 97); -- rb {:board 18, :ch 4} <- ltb {:board 13, :ch 4} ::: {:station "cortina", :ltb-harting 2, :paddle-number 153, :ltb-num+channel {:board 13, :ch 4}, :rb-num+channel {:board 18, :ch 4}, :dsi-slot 3, :panel-number 19, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(196) <= hits_bitmap_i( 98); -- rb {:board 18, :ch 5} <- ltb {:board 13, :ch 5} ::: {:station "cortina", :ltb-harting 2, :paddle-number 154, :ltb-num+channel {:board 13, :ch 5}, :rb-num+channel {:board 18, :ch 5}, :dsi-slot 3, :panel-number 19, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(197) <= hits_bitmap_i( 98); -- rb {:board 18, :ch 6} <- ltb {:board 13, :ch 6} ::: {:station "cortina", :ltb-harting 2, :paddle-number 154, :ltb-num+channel {:board 13, :ch 6}, :rb-num+channel {:board 18, :ch 6}, :dsi-slot 3, :panel-number 19, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(198) <= hits_bitmap_i(102); -- rb {:board 18, :ch 7} <- ltb {:board 13, :ch 13} ::: {:station "cube_corner", :ltb-harting 2, :paddle-number 58, :ltb-num+channel {:board 13, :ch 13}, :rb-num+channel {:board 18, :ch 7}, :dsi-slot 3, :panel-number "E-X135", :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(199) <= hits_bitmap_i(102); -- rb {:board 18, :ch 8} <- ltb {:board 13, :ch 14} ::: {:station "cube_corner", :ltb-harting 2, :paddle-number 58, :ltb-num+channel {:board 13, :ch 14}, :rb-num+channel {:board 18, :ch 8}, :dsi-slot 3, :panel-number "E-X135", :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(200) <= hits_bitmap_i( 99); -- rb {:board 9, :ch 1} <- ltb {:board 13, :ch 7} ::: {:station "cortina", :ltb-harting 2, :paddle-number 133, :ltb-num+channel {:board 13, :ch 7}, :rb-num+channel {:board 9, :ch 1}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(201) <= hits_bitmap_i( 99); -- rb {:board 9, :ch 2} <- ltb {:board 13, :ch 8} ::: {:station "cortina", :ltb-harting 2, :paddle-number 133, :ltb-num+channel {:board 13, :ch 8}, :rb-num+channel {:board 9, :ch 2}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(202) <= hits_bitmap_i(100); -- rb {:board 9, :ch 3} <- ltb {:board 13, :ch 9} ::: {:station "cortina", :ltb-harting 2, :paddle-number 134, :ltb-num+channel {:board 13, :ch 9}, :rb-num+channel {:board 9, :ch 3}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(203) <= hits_bitmap_i(100); -- rb {:board 9, :ch 4} <- ltb {:board 13, :ch 10} ::: {:station "cortina", :ltb-harting 2, :paddle-number 134, :ltb-num+channel {:board 13, :ch 10}, :rb-num+channel {:board 9, :ch 4}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(204) <= hits_bitmap_i(101); -- rb {:board 9, :ch 5} <- ltb {:board 13, :ch 11} ::: {:station "cortina", :ltb-harting 2, :paddle-number 135, :ltb-num+channel {:board 13, :ch 11}, :rb-num+channel {:board 9, :ch 5}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(205) <= hits_bitmap_i(101); -- rb {:board 9, :ch 6} <- ltb {:board 13, :ch 12} ::: {:station "cortina", :ltb-harting 2, :paddle-number 135, :ltb-num+channel {:board 13, :ch 12}, :rb-num+channel {:board 9, :ch 6}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(206) <= hits_bitmap_i(103); -- rb {:board 9, :ch 7} <- ltb {:board 13, :ch 15} ::: {:station "cortina", :ltb-harting 2, :paddle-number 127, :ltb-num+channel {:board 13, :ch 15}, :rb-num+channel {:board 9, :ch 7}, :dsi-slot 3, :panel-number 15, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(207) <= hits_bitmap_i(103); -- rb {:board 9, :ch 8} <- ltb {:board 13, :ch 16} ::: {:station "cortina", :ltb-harting 2, :paddle-number 127, :ltb-num+channel {:board 13, :ch 16}, :rb-num+channel {:board 9, :ch 8}, :dsi-slot 3, :panel-number 15, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(208) <= hits_bitmap_i(105); -- rb {:board 22, :ch 1} <- ltb {:board 14, :ch 3} ::: {:station "cortina", :ltb-harting 3, :paddle-number 132, :ltb-num+channel {:board 14, :ch 3}, :rb-num+channel {:board 22, :ch 1}, :dsi-slot 3, :panel-number 16, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(209) <= hits_bitmap_i(105); -- rb {:board 22, :ch 2} <- ltb {:board 14, :ch 4} ::: {:station "cortina", :ltb-harting 3, :paddle-number 132, :ltb-num+channel {:board 14, :ch 4}, :rb-num+channel {:board 22, :ch 2}, :dsi-slot 3, :panel-number 16, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(210) <= hits_bitmap_i(107); -- rb {:board 22, :ch 3} <- ltb {:board 14, :ch 7} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 20, :ltb-num+channel {:board 14, :ch 7}, :rb-num+channel {:board 22, :ch 3}, :dsi-slot 3, :panel-number 2, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(211) <= hits_bitmap_i(107); -- rb {:board 22, :ch 4} <- ltb {:board 14, :ch 8} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 20, :ltb-num+channel {:board 14, :ch 8}, :rb-num+channel {:board 22, :ch 4}, :dsi-slot 3, :panel-number 2, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(212) <= hits_bitmap_i(109); -- rb {:board 22, :ch 5} <- ltb {:board 14, :ch 11} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 22, :ltb-num+channel {:board 14, :ch 11}, :rb-num+channel {:board 22, :ch 5}, :dsi-slot 3, :panel-number 2, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(213) <= hits_bitmap_i(109); -- rb {:board 22, :ch 6} <- ltb {:board 14, :ch 12} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 22, :ltb-num+channel {:board 14, :ch 12}, :rb-num+channel {:board 22, :ch 6}, :dsi-slot 3, :panel-number 2, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(214) <= hits_bitmap_i(111); -- rb {:board 22, :ch 7} <- ltb {:board 14, :ch 15} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 24, :ltb-num+channel {:board 14, :ch 15}, :rb-num+channel {:board 22, :ch 7}, :dsi-slot 3, :panel-number 2, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(215) <= hits_bitmap_i(111); -- rb {:board 22, :ch 8} <- ltb {:board 14, :ch 16} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 24, :ltb-num+channel {:board 14, :ch 16}, :rb-num+channel {:board 22, :ch 8}, :dsi-slot 3, :panel-number 2, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(216) <= hits_bitmap_i(104); -- rb {:board 26, :ch 1} <- ltb {:board 14, :ch 1} ::: {:station "cortina", :ltb-harting 3, :paddle-number 131, :ltb-num+channel {:board 14, :ch 1}, :rb-num+channel {:board 26, :ch 1}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(217) <= hits_bitmap_i(104); -- rb {:board 26, :ch 2} <- ltb {:board 14, :ch 2} ::: {:station "cortina", :ltb-harting 3, :paddle-number 131, :ltb-num+channel {:board 14, :ch 2}, :rb-num+channel {:board 26, :ch 2}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(218) <= hits_bitmap_i(106); -- rb {:board 26, :ch 3} <- ltb {:board 14, :ch 5} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 19, :ltb-num+channel {:board 14, :ch 5}, :rb-num+channel {:board 26, :ch 3}, :dsi-slot 3, :panel-number 2, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(219) <= hits_bitmap_i(106); -- rb {:board 26, :ch 4} <- ltb {:board 14, :ch 6} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 19, :ltb-num+channel {:board 14, :ch 6}, :rb-num+channel {:board 26, :ch 4}, :dsi-slot 3, :panel-number 2, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(220) <= hits_bitmap_i(108); -- rb {:board 26, :ch 5} <- ltb {:board 14, :ch 9} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 21, :ltb-num+channel {:board 14, :ch 9}, :rb-num+channel {:board 26, :ch 5}, :dsi-slot 3, :panel-number 2, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(221) <= hits_bitmap_i(108); -- rb {:board 26, :ch 6} <- ltb {:board 14, :ch 10} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 21, :ltb-num+channel {:board 14, :ch 10}, :rb-num+channel {:board 26, :ch 6}, :dsi-slot 3, :panel-number 2, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(222) <= hits_bitmap_i(110); -- rb {:board 26, :ch 7} <- ltb {:board 14, :ch 13} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 23, :ltb-num+channel {:board 14, :ch 13}, :rb-num+channel {:board 26, :ch 7}, :dsi-slot 3, :panel-number 2, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(223) <= hits_bitmap_i(110); -- rb {:board 26, :ch 8} <- ltb {:board 14, :ch 14} ::: {:station "cube_bot", :ltb-harting 3, :paddle-number 23, :ltb-num+channel {:board 14, :ch 14}, :rb-num+channel {:board 26, :ch 8}, :dsi-slot 3, :panel-number 2, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(224) <= hits_bitmap_i(113); -- rb {:board 4, :ch 1} <- ltb {:board 15, :ch 3} ::: {:station "cortina", :ltb-harting 4, :paddle-number 130, :ltb-num+channel {:board 15, :ch 3}, :rb-num+channel {:board 4, :ch 1}, :dsi-slot 3, :panel-number 16, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(225) <= hits_bitmap_i(113); -- rb {:board 4, :ch 2} <- ltb {:board 15, :ch 4} ::: {:station "cortina", :ltb-harting 4, :paddle-number 130, :ltb-num+channel {:board 15, :ch 4}, :rb-num+channel {:board 4, :ch 2}, :dsi-slot 3, :panel-number 16, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(226) <= hits_bitmap_i(115); -- rb {:board 4, :ch 3} <- ltb {:board 15, :ch 7} ::: {:station "cube", :ltb-harting 4, :paddle-number 44, :ltb-num+channel {:board 15, :ch 7}, :rb-num+channel {:board 4, :ch 3}, :dsi-slot 3, :panel-number 5, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(227) <= hits_bitmap_i(115); -- rb {:board 4, :ch 4} <- ltb {:board 15, :ch 8} ::: {:station "cube", :ltb-harting 4, :paddle-number 44, :ltb-num+channel {:board 15, :ch 8}, :rb-num+channel {:board 4, :ch 4}, :dsi-slot 3, :panel-number 5, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(228) <= hits_bitmap_i(117); -- rb {:board 4, :ch 5} <- ltb {:board 15, :ch 11} ::: {:station "cube", :ltb-harting 4, :paddle-number 46, :ltb-num+channel {:board 15, :ch 11}, :rb-num+channel {:board 4, :ch 5}, :dsi-slot 3, :panel-number 5, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(229) <= hits_bitmap_i(117); -- rb {:board 4, :ch 6} <- ltb {:board 15, :ch 12} ::: {:station "cube", :ltb-harting 4, :paddle-number 46, :ltb-num+channel {:board 15, :ch 12}, :rb-num+channel {:board 4, :ch 6}, :dsi-slot 3, :panel-number 5, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(230) <= hits_bitmap_i(119); -- rb {:board 4, :ch 7} <- ltb {:board 15, :ch 15} ::: {:station "cube", :ltb-harting 4, :paddle-number 48, :ltb-num+channel {:board 15, :ch 15}, :rb-num+channel {:board 4, :ch 7}, :dsi-slot 3, :panel-number 5, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(231) <= hits_bitmap_i(119); -- rb {:board 4, :ch 8} <- ltb {:board 15, :ch 16} ::: {:station "cube", :ltb-harting 4, :paddle-number 48, :ltb-num+channel {:board 15, :ch 16}, :rb-num+channel {:board 4, :ch 8}, :dsi-slot 3, :panel-number 5, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(232) <= hits_bitmap_i(112); -- rb {:board 2, :ch 1} <- ltb {:board 15, :ch 1} ::: {:station "cortina", :ltb-harting 4, :paddle-number 129, :ltb-num+channel {:board 15, :ch 1}, :rb-num+channel {:board 2, :ch 1}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(233) <= hits_bitmap_i(112); -- rb {:board 2, :ch 2} <- ltb {:board 15, :ch 2} ::: {:station "cortina", :ltb-harting 4, :paddle-number 129, :ltb-num+channel {:board 15, :ch 2}, :rb-num+channel {:board 2, :ch 2}, :dsi-slot 3, :panel-number 16, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(234) <= hits_bitmap_i(114); -- rb {:board 2, :ch 3} <- ltb {:board 15, :ch 5} ::: {:station "cube", :ltb-harting 4, :paddle-number 43, :ltb-num+channel {:board 15, :ch 5}, :rb-num+channel {:board 2, :ch 3}, :dsi-slot 3, :panel-number 5, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(235) <= hits_bitmap_i(114); -- rb {:board 2, :ch 4} <- ltb {:board 15, :ch 6} ::: {:station "cube", :ltb-harting 4, :paddle-number 43, :ltb-num+channel {:board 15, :ch 6}, :rb-num+channel {:board 2, :ch 4}, :dsi-slot 3, :panel-number 5, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(236) <= hits_bitmap_i(116); -- rb {:board 2, :ch 5} <- ltb {:board 15, :ch 9} ::: {:station "cube", :ltb-harting 4, :paddle-number 45, :ltb-num+channel {:board 15, :ch 9}, :rb-num+channel {:board 2, :ch 5}, :dsi-slot 3, :panel-number 5, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(237) <= hits_bitmap_i(116); -- rb {:board 2, :ch 6} <- ltb {:board 15, :ch 10} ::: {:station "cube", :ltb-harting 4, :paddle-number 45, :ltb-num+channel {:board 15, :ch 10}, :rb-num+channel {:board 2, :ch 6}, :dsi-slot 3, :panel-number 5, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(238) <= hits_bitmap_i(118); -- rb {:board 2, :ch 7} <- ltb {:board 15, :ch 13} ::: {:station "cube", :ltb-harting 4, :paddle-number 47, :ltb-num+channel {:board 15, :ch 13}, :rb-num+channel {:board 2, :ch 7}, :dsi-slot 3, :panel-number 5, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(239) <= hits_bitmap_i(118); -- rb {:board 2, :ch 8} <- ltb {:board 15, :ch 14} ::: {:station "cube", :ltb-harting 4, :paddle-number 47, :ltb-num+channel {:board 15, :ch 14}, :rb-num+channel {:board 2, :ch 8}, :dsi-slot 3, :panel-number 5, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(240) <= hits_bitmap_i(120); -- rb {:board 44, :ch 1} <- ltb {:board 16, :ch 1} ::: {:station "cube", :ltb-harting 0, :paddle-number 42, :ltb-num+channel {:board 16, :ch 1}, :rb-num+channel {:board 44, :ch 1}, :dsi-slot 4, :panel-number 5, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(241) <= hits_bitmap_i(120); -- rb {:board 44, :ch 2} <- ltb {:board 16, :ch 2} ::: {:station "cube", :ltb-harting 0, :paddle-number 42, :ltb-num+channel {:board 16, :ch 2}, :rb-num+channel {:board 44, :ch 2}, :dsi-slot 4, :panel-number 5, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(242) <= hits_bitmap_i(122); -- rb {:board 44, :ch 3} <- ltb {:board 16, :ch 5} ::: {:station "cube", :ltb-harting 0, :paddle-number 12, :ltb-num+channel {:board 16, :ch 5}, :rb-num+channel {:board 44, :ch 3}, :dsi-slot 4, :panel-number 1, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(243) <= hits_bitmap_i(122); -- rb {:board 44, :ch 4} <- ltb {:board 16, :ch 6} ::: {:station "cube", :ltb-harting 0, :paddle-number 12, :ltb-num+channel {:board 16, :ch 6}, :rb-num+channel {:board 44, :ch 4}, :dsi-slot 4, :panel-number 1, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(244) <= hits_bitmap_i(124); -- rb {:board 44, :ch 5} <- ltb {:board 16, :ch 9} ::: {:station "cube", :ltb-harting 0, :paddle-number 10, :ltb-num+channel {:board 16, :ch 9}, :rb-num+channel {:board 44, :ch 5}, :dsi-slot 4, :panel-number 1, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(245) <= hits_bitmap_i(124); -- rb {:board 44, :ch 6} <- ltb {:board 16, :ch 10} ::: {:station "cube", :ltb-harting 0, :paddle-number 10, :ltb-num+channel {:board 16, :ch 10}, :rb-num+channel {:board 44, :ch 6}, :dsi-slot 4, :panel-number 1, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(246) <= hits_bitmap_i(126); -- rb {:board 44, :ch 7} <- ltb {:board 16, :ch 13} ::: {:station "cube", :ltb-harting 0, :paddle-number 8, :ltb-num+channel {:board 16, :ch 13}, :rb-num+channel {:board 44, :ch 7}, :dsi-slot 4, :panel-number 1, :harting-half :A, :paddle-end :B, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(247) <= hits_bitmap_i(126); -- rb {:board 44, :ch 8} <- ltb {:board 16, :ch 14} ::: {:station "cube", :ltb-harting 0, :paddle-number 8, :ltb-num+channel {:board 16, :ch 14}, :rb-num+channel {:board 44, :ch 8}, :dsi-slot 4, :panel-number 1, :harting-half :A, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(248) <= hits_bitmap_i(121); -- rb {:board 30, :ch 1} <- ltb {:board 16, :ch 3} ::: {:station "cube", :ltb-harting 0, :paddle-number 41, :ltb-num+channel {:board 16, :ch 3}, :rb-num+channel {:board 30, :ch 1}, :dsi-slot 4, :panel-number 5, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(249) <= hits_bitmap_i(121); -- rb {:board 30, :ch 2} <- ltb {:board 16, :ch 4} ::: {:station "cube", :ltb-harting 0, :paddle-number 41, :ltb-num+channel {:board 16, :ch 4}, :rb-num+channel {:board 30, :ch 2}, :dsi-slot 4, :panel-number 5, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(250) <= hits_bitmap_i(123); -- rb {:board 30, :ch 3} <- ltb {:board 16, :ch 7} ::: {:station "cube", :ltb-harting 0, :paddle-number 11, :ltb-num+channel {:board 16, :ch 7}, :rb-num+channel {:board 30, :ch 3}, :dsi-slot 4, :panel-number 1, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(251) <= hits_bitmap_i(123); -- rb {:board 30, :ch 4} <- ltb {:board 16, :ch 8} ::: {:station "cube", :ltb-harting 0, :paddle-number 11, :ltb-num+channel {:board 16, :ch 8}, :rb-num+channel {:board 30, :ch 4}, :dsi-slot 4, :panel-number 1, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(252) <= hits_bitmap_i(125); -- rb {:board 30, :ch 5} <- ltb {:board 16, :ch 11} ::: {:station "cube", :ltb-harting 0, :paddle-number 9, :ltb-num+channel {:board 16, :ch 11}, :rb-num+channel {:board 30, :ch 5}, :dsi-slot 4, :panel-number 1, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(253) <= hits_bitmap_i(125); -- rb {:board 30, :ch 6} <- ltb {:board 16, :ch 12} ::: {:station "cube", :ltb-harting 0, :paddle-number 9, :ltb-num+channel {:board 16, :ch 12}, :rb-num+channel {:board 30, :ch 6}, :dsi-slot 4, :panel-number 1, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(254) <= hits_bitmap_i(127); -- rb {:board 30, :ch 7} <- ltb {:board 16, :ch 15} ::: {:station "cube", :ltb-harting 0, :paddle-number 7, :ltb-num+channel {:board 16, :ch 15}, :rb-num+channel {:board 30, :ch 7}, :dsi-slot 4, :panel-number 1, :harting-half :B, :paddle-end :B, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(255) <= hits_bitmap_i(127); -- rb {:board 30, :ch 8} <- ltb {:board 16, :ch 16} ::: {:station "cube", :ltb-harting 0, :paddle-number 7, :ltb-num+channel {:board 16, :ch 16}, :rb-num+channel {:board 30, :ch 8}, :dsi-slot 4, :panel-number 1, :harting-half :B, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(256) <= hits_bitmap_i(129); -- rb {:board 17, :ch 1} <- ltb {:board 17, :ch 3} ::: {:station "cube_corner", :ltb-harting 1, :paddle-number 59, :ltb-num+channel {:board 17, :ch 3}, :rb-num+channel {:board 17, :ch 1}, :dsi-slot 4, :panel-number "E-X225", :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(257) <= hits_bitmap_i(129); -- rb {:board 17, :ch 2} <- ltb {:board 17, :ch 4} ::: {:station "cube_corner", :ltb-harting 1, :paddle-number 59, :ltb-num+channel {:board 17, :ch 4}, :rb-num+channel {:board 17, :ch 2}, :dsi-slot 4, :panel-number "E-X225", :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(258) <= hits_bitmap_i(130); -- rb {:board 17, :ch 3} <- ltb {:board 17, :ch 5} ::: {:station "cortina", :ltb-harting 1, :paddle-number 155, :ltb-num+channel {:board 17, :ch 5}, :rb-num+channel {:board 17, :ch 3}, :dsi-slot 4, :panel-number 20, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(259) <= hits_bitmap_i(135); -- rb {:board 17, :ch 4} <- ltb {:board 17, :ch 16} ::: {:station "cortina", :ltb-harting 1, :paddle-number 155, :ltb-num+channel {:board 17, :ch 16}, :rb-num+channel {:board 17, :ch 4}, :dsi-slot 4, :panel-number 20, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(260) <= hits_bitmap_i(132); -- rb {:board 17, :ch 5} <- ltb {:board 17, :ch 9} ::: {:station "cortina", :ltb-harting 1, :paddle-number 157, :ltb-num+channel {:board 17, :ch 9}, :rb-num+channel {:board 17, :ch 5}, :dsi-slot 4, :panel-number 20, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(261) <= hits_bitmap_i(132); -- rb {:board 17, :ch 6} <- ltb {:board 17, :ch 10} ::: {:station "cortina", :ltb-harting 1, :paddle-number 157, :ltb-num+channel {:board 17, :ch 10}, :rb-num+channel {:board 17, :ch 6}, :dsi-slot 4, :panel-number 20, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(262) <= hits_bitmap_i(134); -- rb {:board 17, :ch 7} <- ltb {:board 17, :ch 13} ::: {:station "cortina", :ltb-harting 1, :paddle-number 137, :ltb-num+channel {:board 17, :ch 13}, :rb-num+channel {:board 17, :ch 7}, :dsi-slot 4, :panel-number 16, :harting-half :A, :paddle-end :B, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(263) <= hits_bitmap_i(134); -- rb {:board 17, :ch 8} <- ltb {:board 17, :ch 14} ::: {:station "cortina", :ltb-harting 1, :paddle-number 137, :ltb-num+channel {:board 17, :ch 14}, :rb-num+channel {:board 17, :ch 8}, :dsi-slot 4, :panel-number 16, :harting-half :A, :paddle-end :A, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(264) <= hits_bitmap_i(128); -- rb {:board 7, :ch 1} <- ltb {:board 17, :ch 1} ::: {:station "cortina", :ltb-harting 1, :paddle-number 147, :ltb-num+channel {:board 17, :ch 1}, :rb-num+channel {:board 7, :ch 1}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(265) <= hits_bitmap_i(128); -- rb {:board 7, :ch 2} <- ltb {:board 17, :ch 2} ::: {:station "cortina", :ltb-harting 1, :paddle-number 147, :ltb-num+channel {:board 17, :ch 2}, :rb-num+channel {:board 7, :ch 2}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(266) <= hits_bitmap_i(131); -- rb {:board 7, :ch 3} <- ltb {:board 17, :ch 7} ::: {:station "cortina", :ltb-harting 1, :paddle-number 156, :ltb-num+channel {:board 17, :ch 7}, :rb-num+channel {:board 7, :ch 3}, :dsi-slot 4, :panel-number 20, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(267) <= hits_bitmap_i(131); -- rb {:board 7, :ch 4} <- ltb {:board 17, :ch 8} ::: {:station "cortina", :ltb-harting 1, :paddle-number 156, :ltb-num+channel {:board 17, :ch 8}, :rb-num+channel {:board 7, :ch 4}, :dsi-slot 4, :panel-number 20, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(268) <= hits_bitmap_i(133); -- rb {:board 7, :ch 5} <- ltb {:board 17, :ch 11} ::: {:station "cortina", :ltb-harting 1, :paddle-number 138, :ltb-num+channel {:board 17, :ch 11}, :rb-num+channel {:board 7, :ch 5}, :dsi-slot 4, :panel-number 16, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(269) <= hits_bitmap_i(133); -- rb {:board 7, :ch 6} <- ltb {:board 17, :ch 12} ::: {:station "cortina", :ltb-harting 1, :paddle-number 138, :ltb-num+channel {:board 17, :ch 12}, :rb-num+channel {:board 7, :ch 6}, :dsi-slot 4, :panel-number 16, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(270) <= hits_bitmap_i(135); -- rb {:board 7, :ch 7} <- ltb {:board 17, :ch 15} ::: {:station "cortina", :ltb-harting 1, :paddle-number 136, :ltb-num+channel {:board 17, :ch 15}, :rb-num+channel {:board 7, :ch 7}, :dsi-slot 4, :panel-number 16, :harting-half :B, :paddle-end :B, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(271) <= hits_bitmap_i(135); -- rb {:board 7, :ch 8} <- ltb {:board 17, :ch 16} ::: {:station "cortina", :ltb-harting 1, :paddle-number 136, :ltb-num+channel {:board 17, :ch 16}, :rb-num+channel {:board 7, :ch 8}, :dsi-slot 4, :panel-number 16, :harting-half :B, :paddle-end :A, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(272) <= hits_bitmap_i(137); -- rb {:board 34, :ch 1} <- ltb {:board 18, :ch 3} ::: {:station "cortina", :ltb-harting 2, :paddle-number 140, :ltb-num+channel {:board 18, :ch 3}, :rb-num+channel {:board 34, :ch 1}, :dsi-slot 4, :panel-number 17, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(273) <= hits_bitmap_i(137); -- rb {:board 34, :ch 2} <- ltb {:board 18, :ch 4} ::: {:station "cortina", :ltb-harting 2, :paddle-number 140, :ltb-num+channel {:board 18, :ch 4}, :rb-num+channel {:board 34, :ch 2}, :dsi-slot 4, :panel-number 17, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(274) <= hits_bitmap_i(139); -- rb {:board 34, :ch 3} <- ltb {:board 18, :ch 7} ::: {:station "cortina", :ltb-harting 2, :paddle-number 142, :ltb-num+channel {:board 18, :ch 7}, :rb-num+channel {:board 34, :ch 3}, :dsi-slot 4, :panel-number 17, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(275) <= hits_bitmap_i(139); -- rb {:board 34, :ch 4} <- ltb {:board 18, :ch 8} ::: {:station "cortina", :ltb-harting 2, :paddle-number 142, :ltb-num+channel {:board 18, :ch 8}, :rb-num+channel {:board 34, :ch 4}, :dsi-slot 4, :panel-number 17, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(276) <= hits_bitmap_i(141); -- rb {:board 34, :ch 5} <- ltb {:board 18, :ch 11} ::: {:station "cortina", :ltb-harting 2, :paddle-number 144, :ltb-num+channel {:board 18, :ch 11}, :rb-num+channel {:board 34, :ch 5}, :dsi-slot 4, :panel-number 17, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(277) <= hits_bitmap_i(141); -- rb {:board 34, :ch 6} <- ltb {:board 18, :ch 12} ::: {:station "cortina", :ltb-harting 2, :paddle-number 144, :ltb-num+channel {:board 18, :ch 12}, :rb-num+channel {:board 34, :ch 6}, :dsi-slot 4, :panel-number 17, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(278) <= hits_bitmap_i(143); -- rb {:board 34, :ch 7} <- ltb {:board 18, :ch 15} ::: {:station "cortina", :ltb-harting 2, :paddle-number 146, :ltb-num+channel {:board 18, :ch 15}, :rb-num+channel {:board 34, :ch 7}, :dsi-slot 4, :panel-number 17, :harting-half :A, :paddle-end :B, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(279) <= hits_bitmap_i(143); -- rb {:board 34, :ch 8} <- ltb {:board 18, :ch 16} ::: {:station "cortina", :ltb-harting 2, :paddle-number 146, :ltb-num+channel {:board 18, :ch 16}, :rb-num+channel {:board 34, :ch 8}, :dsi-slot 4, :panel-number 17, :harting-half :A, :paddle-end :A, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(280) <= hits_bitmap_i(136); -- rb {:board 33, :ch 1} <- ltb {:board 18, :ch 1} ::: {:station "cortina", :ltb-harting 2, :paddle-number 139, :ltb-num+channel {:board 18, :ch 1}, :rb-num+channel {:board 33, :ch 1}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(281) <= hits_bitmap_i(136); -- rb {:board 33, :ch 2} <- ltb {:board 18, :ch 2} ::: {:station "cortina", :ltb-harting 2, :paddle-number 139, :ltb-num+channel {:board 18, :ch 2}, :rb-num+channel {:board 33, :ch 2}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(282) <= hits_bitmap_i(138); -- rb {:board 33, :ch 3} <- ltb {:board 18, :ch 5} ::: {:station "cortina", :ltb-harting 2, :paddle-number 141, :ltb-num+channel {:board 18, :ch 5}, :rb-num+channel {:board 33, :ch 3}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(283) <= hits_bitmap_i(138); -- rb {:board 33, :ch 4} <- ltb {:board 18, :ch 6} ::: {:station "cortina", :ltb-harting 2, :paddle-number 141, :ltb-num+channel {:board 18, :ch 6}, :rb-num+channel {:board 33, :ch 4}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(284) <= hits_bitmap_i(140); -- rb {:board 33, :ch 5} <- ltb {:board 18, :ch 9} ::: {:station "cortina", :ltb-harting 2, :paddle-number 143, :ltb-num+channel {:board 18, :ch 9}, :rb-num+channel {:board 33, :ch 5}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(285) <= hits_bitmap_i(140); -- rb {:board 33, :ch 6} <- ltb {:board 18, :ch 10} ::: {:station "cortina", :ltb-harting 2, :paddle-number 143, :ltb-num+channel {:board 18, :ch 10}, :rb-num+channel {:board 33, :ch 6}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(286) <= hits_bitmap_i(142); -- rb {:board 33, :ch 7} <- ltb {:board 18, :ch 13} ::: {:station "cortina", :ltb-harting 2, :paddle-number 145, :ltb-num+channel {:board 18, :ch 13}, :rb-num+channel {:board 33, :ch 7}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :B, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(287) <= hits_bitmap_i(142); -- rb {:board 33, :ch 8} <- ltb {:board 18, :ch 14} ::: {:station "cortina", :ltb-harting 2, :paddle-number 145, :ltb-num+channel {:board 18, :ch 14}, :rb-num+channel {:board 33, :ch 8}, :dsi-slot 4, :panel-number 17, :harting-half :B, :paddle-end :A, :rb-harting 2, :rat-number 18}
  rb_ch_bitmap_o(288) <= hits_bitmap_i(144); -- rb {:board 6, :ch 1} <- ltb {:board 19, :ch 1} ::: {:station "cube", :ltb-harting 3, :paddle-number 56, :ltb-num+channel {:board 19, :ch 1}, :rb-num+channel {:board 6, :ch 1}, :dsi-slot 4, :panel-number 6, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(289) <= hits_bitmap_i(144); -- rb {:board 6, :ch 2} <- ltb {:board 19, :ch 2} ::: {:station "cube", :ltb-harting 3, :paddle-number 56, :ltb-num+channel {:board 19, :ch 2}, :rb-num+channel {:board 6, :ch 2}, :dsi-slot 4, :panel-number 6, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(290) <= hits_bitmap_i(145); -- rb {:board 6, :ch 3} <- ltb {:board 19, :ch 3} ::: {:station "cube", :ltb-harting 3, :paddle-number 54, :ltb-num+channel {:board 19, :ch 3}, :rb-num+channel {:board 6, :ch 3}, :dsi-slot 4, :panel-number 6, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(291) <= hits_bitmap_i(145); -- rb {:board 6, :ch 4} <- ltb {:board 19, :ch 4} ::: {:station "cube", :ltb-harting 3, :paddle-number 54, :ltb-num+channel {:board 19, :ch 4}, :rb-num+channel {:board 6, :ch 4}, :dsi-slot 4, :panel-number 6, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(292) <= hits_bitmap_i(146); -- rb {:board 6, :ch 5} <- ltb {:board 19, :ch 5} ::: {:station "cube", :ltb-harting 3, :paddle-number 52, :ltb-num+channel {:board 19, :ch 5}, :rb-num+channel {:board 6, :ch 5}, :dsi-slot 4, :panel-number 6, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(293) <= hits_bitmap_i(146); -- rb {:board 6, :ch 6} <- ltb {:board 19, :ch 6} ::: {:station "cube", :ltb-harting 3, :paddle-number 52, :ltb-num+channel {:board 19, :ch 6}, :rb-num+channel {:board 6, :ch 6}, :dsi-slot 4, :panel-number 6, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(294) <= hits_bitmap_i(147); -- rb {:board 6, :ch 7} <- ltb {:board 19, :ch 7} ::: {:station "cube", :ltb-harting 3, :paddle-number 50, :ltb-num+channel {:board 19, :ch 7}, :rb-num+channel {:board 6, :ch 7}, :dsi-slot 4, :panel-number 6, :harting-half :A, :paddle-end :B, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(295) <= hits_bitmap_i(147); -- rb {:board 6, :ch 8} <- ltb {:board 19, :ch 8} ::: {:station "cube", :ltb-harting 3, :paddle-number 50, :ltb-num+channel {:board 19, :ch 8}, :rb-num+channel {:board 6, :ch 8}, :dsi-slot 4, :panel-number 6, :harting-half :A, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(296) <= hits_bitmap_i(151); -- rb {:board 36, :ch 1} <- ltb {:board 19, :ch 15} ::: {:station "cube", :ltb-harting 3, :paddle-number 55, :ltb-num+channel {:board 19, :ch 15}, :rb-num+channel {:board 36, :ch 1}, :dsi-slot 4, :panel-number 6, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(297) <= hits_bitmap_i(151); -- rb {:board 36, :ch 2} <- ltb {:board 19, :ch 16} ::: {:station "cube", :ltb-harting 3, :paddle-number 55, :ltb-num+channel {:board 19, :ch 16}, :rb-num+channel {:board 36, :ch 2}, :dsi-slot 4, :panel-number 6, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(298) <= hits_bitmap_i(150); -- rb {:board 36, :ch 3} <- ltb {:board 19, :ch 13} ::: {:station "cube", :ltb-harting 3, :paddle-number 53, :ltb-num+channel {:board 19, :ch 13}, :rb-num+channel {:board 36, :ch 3}, :dsi-slot 4, :panel-number 6, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(299) <= hits_bitmap_i(150); -- rb {:board 36, :ch 4} <- ltb {:board 19, :ch 14} ::: {:station "cube", :ltb-harting 3, :paddle-number 53, :ltb-num+channel {:board 19, :ch 14}, :rb-num+channel {:board 36, :ch 4}, :dsi-slot 4, :panel-number 6, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(300) <= hits_bitmap_i(149); -- rb {:board 36, :ch 5} <- ltb {:board 19, :ch 11} ::: {:station "cube", :ltb-harting 3, :paddle-number 51, :ltb-num+channel {:board 19, :ch 11}, :rb-num+channel {:board 36, :ch 5}, :dsi-slot 4, :panel-number 6, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(301) <= hits_bitmap_i(149); -- rb {:board 36, :ch 6} <- ltb {:board 19, :ch 12} ::: {:station "cube", :ltb-harting 3, :paddle-number 51, :ltb-num+channel {:board 19, :ch 12}, :rb-num+channel {:board 36, :ch 6}, :dsi-slot 4, :panel-number 6, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(302) <= hits_bitmap_i(148); -- rb {:board 36, :ch 7} <- ltb {:board 19, :ch 9} ::: {:station "cube", :ltb-harting 3, :paddle-number 49, :ltb-num+channel {:board 19, :ch 9}, :rb-num+channel {:board 36, :ch 7}, :dsi-slot 4, :panel-number 6, :harting-half :B, :paddle-end :B, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(303) <= hits_bitmap_i(148); -- rb {:board 36, :ch 8} <- ltb {:board 19, :ch 10} ::: {:station "cube", :ltb-harting 3, :paddle-number 49, :ltb-num+channel {:board 19, :ch 10}, :rb-num+channel {:board 36, :ch 8}, :dsi-slot 4, :panel-number 6, :harting-half :B, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(304) <= hits_bitmap_i(152); -- rb {:board 5, :ch 1} <- ltb {:board 20, :ch 1} ::: {:station "cortina", :ltb-harting 4, :paddle-number 126, :ltb-num+channel {:board 20, :ch 1}, :rb-num+channel {:board 5, :ch 1}, :dsi-slot 4, :panel-number 15, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(305) <= hits_bitmap_i(152); -- rb {:board 5, :ch 2} <- ltb {:board 20, :ch 2} ::: {:station "cortina", :ltb-harting 4, :paddle-number 126, :ltb-num+channel {:board 20, :ch 2}, :rb-num+channel {:board 5, :ch 2}, :dsi-slot 4, :panel-number 15, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(306) <= hits_bitmap_i(154); -- rb {:board 5, :ch 3} <- ltb {:board 20, :ch 5} ::: {:station "cortina", :ltb-harting 4, :paddle-number 124, :ltb-num+channel {:board 20, :ch 5}, :rb-num+channel {:board 5, :ch 3}, :dsi-slot 4, :panel-number 15, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(307) <= hits_bitmap_i(154); -- rb {:board 5, :ch 4} <- ltb {:board 20, :ch 6} ::: {:station "cortina", :ltb-harting 4, :paddle-number 124, :ltb-num+channel {:board 20, :ch 6}, :rb-num+channel {:board 5, :ch 4}, :dsi-slot 4, :panel-number 15, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(308) <= hits_bitmap_i(156); -- rb {:board 5, :ch 5} <- ltb {:board 20, :ch 9} ::: {:station "cortina", :ltb-harting 4, :paddle-number 122, :ltb-num+channel {:board 20, :ch 9}, :rb-num+channel {:board 5, :ch 5}, :dsi-slot 4, :panel-number 15, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(309) <= hits_bitmap_i(156); -- rb {:board 5, :ch 6} <- ltb {:board 20, :ch 10} ::: {:station "cortina", :ltb-harting 4, :paddle-number 122, :ltb-num+channel {:board 20, :ch 10}, :rb-num+channel {:board 5, :ch 6}, :dsi-slot 4, :panel-number 15, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(310) <= hits_bitmap_i(158); -- rb {:board 5, :ch 7} <- ltb {:board 20, :ch 13} ::: {:station "cortina", :ltb-harting 4, :paddle-number 120, :ltb-num+channel {:board 20, :ch 13}, :rb-num+channel {:board 5, :ch 7}, :dsi-slot 4, :panel-number 15, :harting-half :A, :paddle-end :B, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(311) <= hits_bitmap_i(158); -- rb {:board 5, :ch 8} <- ltb {:board 20, :ch 14} ::: {:station "cortina", :ltb-harting 4, :paddle-number 120, :ltb-num+channel {:board 20, :ch 14}, :rb-num+channel {:board 5, :ch 8}, :dsi-slot 4, :panel-number 15, :harting-half :A, :paddle-end :A, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(312) <= hits_bitmap_i(153); -- rb {:board 28, :ch 1} <- ltb {:board 20, :ch 3} ::: {:station "cortina", :ltb-harting 4, :paddle-number 125, :ltb-num+channel {:board 20, :ch 3}, :rb-num+channel {:board 28, :ch 1}, :dsi-slot 4, :panel-number 15, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(313) <= hits_bitmap_i(153); -- rb {:board 28, :ch 2} <- ltb {:board 20, :ch 4} ::: {:station "cortina", :ltb-harting 4, :paddle-number 125, :ltb-num+channel {:board 20, :ch 4}, :rb-num+channel {:board 28, :ch 2}, :dsi-slot 4, :panel-number 15, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(314) <= hits_bitmap_i(155); -- rb {:board 28, :ch 3} <- ltb {:board 20, :ch 7} ::: {:station "cortina", :ltb-harting 4, :paddle-number 123, :ltb-num+channel {:board 20, :ch 7}, :rb-num+channel {:board 28, :ch 3}, :dsi-slot 4, :panel-number 15, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(315) <= hits_bitmap_i(155); -- rb {:board 28, :ch 4} <- ltb {:board 20, :ch 8} ::: {:station "cortina", :ltb-harting 4, :paddle-number 123, :ltb-num+channel {:board 20, :ch 8}, :rb-num+channel {:board 28, :ch 4}, :dsi-slot 4, :panel-number 15, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(316) <= hits_bitmap_i(157); -- rb {:board 28, :ch 5} <- ltb {:board 20, :ch 11} ::: {:station "cortina", :ltb-harting 4, :paddle-number 121, :ltb-num+channel {:board 20, :ch 11}, :rb-num+channel {:board 28, :ch 5}, :dsi-slot 4, :panel-number 15, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(317) <= hits_bitmap_i(157); -- rb {:board 28, :ch 6} <- ltb {:board 20, :ch 12} ::: {:station "cortina", :ltb-harting 4, :paddle-number 121, :ltb-num+channel {:board 20, :ch 12}, :rb-num+channel {:board 28, :ch 6}, :dsi-slot 4, :panel-number 15, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(318) <= hits_bitmap_i(159); -- rb {:board 28, :ch 7} <- ltb {:board 20, :ch 15} ::: {:station "cortina", :ltb-harting 4, :paddle-number 119, :ltb-num+channel {:board 20, :ch 15}, :rb-num+channel {:board 28, :ch 7}, :dsi-slot 4, :panel-number 15, :harting-half :B, :paddle-end :B, :rb-harting 4, :rat-number 20}
  rb_ch_bitmap_o(319) <= hits_bitmap_i(159); -- rb {:board 28, :ch 8} <- ltb {:board 20, :ch 16} ::: {:station "cortina", :ltb-harting 4, :paddle-number 119, :ltb-num+channel {:board 20, :ch 16}, :rb-num+channel {:board 28, :ch 8}, :dsi-slot 4, :panel-number 15, :harting-half :B, :paddle-end :A, :rb-harting 4, :rat-number 20}
  --END: autoinsert mapping

end behavioral;
