library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.types_pkg.all;
use work.mt_types.all;
use work.constants.all;
use work.components.all;

-- Panel mapping: https://docs.google.com/spreadsheets/d/1i41fsmLf7IjfYbr1coTo9V4uk3t1GXAGgt0aOeCkeeA/edit#gid=0

entity trigger_top is
  generic (DEBUG : boolean := true);
  port(


    clk : in std_logic;

    reset : in std_logic;

    event_cnt_reset : in std_logic;

    any_hit_trigger_is_global : in std_logic;
    track_trigger_is_global   : in std_logic;
    track_central_is_global   : in std_logic;

    any_hit_trigger_prescale : in std_logic_vector (31 downto 0);
    track_trigger_prescale   : in std_logic_vector (31 downto 0);
    track_central_prescale   : in std_logic_vector (31 downto 0);

    hit_thresh : in std_logic_vector (1 downto 0);

    read_all_channels : in std_logic := '1';

    -- this is an array of 25*8 = 200 thresholds, where each threshold is a 2
    -- bit value
    hits_i_0 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_1 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_2 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_3 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_4 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_5 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_6 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_7 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_8 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_9 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_10 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_11 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_12 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_13 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_14 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_15 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_16 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_17 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_18 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_19 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_20 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_21 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_22 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_23 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_24 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_25 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_26 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_27 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_28 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_29 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_30 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_31 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_32 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_33 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_34 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_35 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_36 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_37 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_38 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_39 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_40 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_41 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_42 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_43 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_44 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_45 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_46 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_47 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_48 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_49 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_50 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_51 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_52 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_53 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_54 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_55 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_56 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_57 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_58 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_59 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_60 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_61 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_62 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_63 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_64 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_65 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_66 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_67 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_68 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_69 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_70 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_71 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_72 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_73 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_74 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_75 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_76 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_77 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_78 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_79 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_80 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_81 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_82 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_83 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_84 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_85 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_86 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_87 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_88 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_89 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_90 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_91 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_92 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_93 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_94 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_95 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_96 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_97 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_98 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_99 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_100 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_101 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_102 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_103 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_104 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_105 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_106 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_107 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_108 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_109 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_110 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_111 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_112 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_113 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_114 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_115 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_116 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_117 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_118 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_119 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_120 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_121 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_122 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_123 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_124 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_125 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_126 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_127 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_128 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_129 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_130 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_131 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_132 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_133 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_134 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_135 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_136 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_137 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_138 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_139 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_140 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_141 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_142 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_143 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_144 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_145 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_146 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_147 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_148 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_149 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_150 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_151 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_152 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_153 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_154 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_155 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_156 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_157 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_158 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_159 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_160 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_161 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_162 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_163 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_164 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_165 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_166 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_167 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_168 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_169 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_170 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_171 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_172 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_173 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_174 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_175 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_176 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_177 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_178 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_179 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_180 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_181 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_182 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_183 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_184 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_185 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_186 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_187 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_188 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_189 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_190 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_191 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_192 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_193 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_194 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_195 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_196 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_197 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_198 : in std_logic_vector(1 downto 0) := (others => '0');
    hits_i_199 : in std_logic_vector(1 downto 0) := (others => '0');

    hits_o_0 : out std_logic_vector(1 downto 0);
    hits_o_1 : out std_logic_vector(1 downto 0);
    hits_o_2 : out std_logic_vector(1 downto 0);
    hits_o_3 : out std_logic_vector(1 downto 0);
    hits_o_4 : out std_logic_vector(1 downto 0);
    hits_o_5 : out std_logic_vector(1 downto 0);
    hits_o_6 : out std_logic_vector(1 downto 0);
    hits_o_7 : out std_logic_vector(1 downto 0);
    hits_o_8 : out std_logic_vector(1 downto 0);
    hits_o_9 : out std_logic_vector(1 downto 0);
    hits_o_10 : out std_logic_vector(1 downto 0);
    hits_o_11 : out std_logic_vector(1 downto 0);
    hits_o_12 : out std_logic_vector(1 downto 0);
    hits_o_13 : out std_logic_vector(1 downto 0);
    hits_o_14 : out std_logic_vector(1 downto 0);
    hits_o_15 : out std_logic_vector(1 downto 0);
    hits_o_16 : out std_logic_vector(1 downto 0);
    hits_o_17 : out std_logic_vector(1 downto 0);
    hits_o_18 : out std_logic_vector(1 downto 0);
    hits_o_19 : out std_logic_vector(1 downto 0);
    hits_o_20 : out std_logic_vector(1 downto 0);
    hits_o_21 : out std_logic_vector(1 downto 0);
    hits_o_22 : out std_logic_vector(1 downto 0);
    hits_o_23 : out std_logic_vector(1 downto 0);
    hits_o_24 : out std_logic_vector(1 downto 0);
    hits_o_25 : out std_logic_vector(1 downto 0);
    hits_o_26 : out std_logic_vector(1 downto 0);
    hits_o_27 : out std_logic_vector(1 downto 0);
    hits_o_28 : out std_logic_vector(1 downto 0);
    hits_o_29 : out std_logic_vector(1 downto 0);
    hits_o_30 : out std_logic_vector(1 downto 0);
    hits_o_31 : out std_logic_vector(1 downto 0);
    hits_o_32 : out std_logic_vector(1 downto 0);
    hits_o_33 : out std_logic_vector(1 downto 0);
    hits_o_34 : out std_logic_vector(1 downto 0);
    hits_o_35 : out std_logic_vector(1 downto 0);
    hits_o_36 : out std_logic_vector(1 downto 0);
    hits_o_37 : out std_logic_vector(1 downto 0);
    hits_o_38 : out std_logic_vector(1 downto 0);
    hits_o_39 : out std_logic_vector(1 downto 0);
    hits_o_40 : out std_logic_vector(1 downto 0);
    hits_o_41 : out std_logic_vector(1 downto 0);
    hits_o_42 : out std_logic_vector(1 downto 0);
    hits_o_43 : out std_logic_vector(1 downto 0);
    hits_o_44 : out std_logic_vector(1 downto 0);
    hits_o_45 : out std_logic_vector(1 downto 0);
    hits_o_46 : out std_logic_vector(1 downto 0);
    hits_o_47 : out std_logic_vector(1 downto 0);
    hits_o_48 : out std_logic_vector(1 downto 0);
    hits_o_49 : out std_logic_vector(1 downto 0);
    hits_o_50 : out std_logic_vector(1 downto 0);
    hits_o_51 : out std_logic_vector(1 downto 0);
    hits_o_52 : out std_logic_vector(1 downto 0);
    hits_o_53 : out std_logic_vector(1 downto 0);
    hits_o_54 : out std_logic_vector(1 downto 0);
    hits_o_55 : out std_logic_vector(1 downto 0);
    hits_o_56 : out std_logic_vector(1 downto 0);
    hits_o_57 : out std_logic_vector(1 downto 0);
    hits_o_58 : out std_logic_vector(1 downto 0);
    hits_o_59 : out std_logic_vector(1 downto 0);
    hits_o_60 : out std_logic_vector(1 downto 0);
    hits_o_61 : out std_logic_vector(1 downto 0);
    hits_o_62 : out std_logic_vector(1 downto 0);
    hits_o_63 : out std_logic_vector(1 downto 0);
    hits_o_64 : out std_logic_vector(1 downto 0);
    hits_o_65 : out std_logic_vector(1 downto 0);
    hits_o_66 : out std_logic_vector(1 downto 0);
    hits_o_67 : out std_logic_vector(1 downto 0);
    hits_o_68 : out std_logic_vector(1 downto 0);
    hits_o_69 : out std_logic_vector(1 downto 0);
    hits_o_70 : out std_logic_vector(1 downto 0);
    hits_o_71 : out std_logic_vector(1 downto 0);
    hits_o_72 : out std_logic_vector(1 downto 0);
    hits_o_73 : out std_logic_vector(1 downto 0);
    hits_o_74 : out std_logic_vector(1 downto 0);
    hits_o_75 : out std_logic_vector(1 downto 0);
    hits_o_76 : out std_logic_vector(1 downto 0);
    hits_o_77 : out std_logic_vector(1 downto 0);
    hits_o_78 : out std_logic_vector(1 downto 0);
    hits_o_79 : out std_logic_vector(1 downto 0);
    hits_o_80 : out std_logic_vector(1 downto 0);
    hits_o_81 : out std_logic_vector(1 downto 0);
    hits_o_82 : out std_logic_vector(1 downto 0);
    hits_o_83 : out std_logic_vector(1 downto 0);
    hits_o_84 : out std_logic_vector(1 downto 0);
    hits_o_85 : out std_logic_vector(1 downto 0);
    hits_o_86 : out std_logic_vector(1 downto 0);
    hits_o_87 : out std_logic_vector(1 downto 0);
    hits_o_88 : out std_logic_vector(1 downto 0);
    hits_o_89 : out std_logic_vector(1 downto 0);
    hits_o_90 : out std_logic_vector(1 downto 0);
    hits_o_91 : out std_logic_vector(1 downto 0);
    hits_o_92 : out std_logic_vector(1 downto 0);
    hits_o_93 : out std_logic_vector(1 downto 0);
    hits_o_94 : out std_logic_vector(1 downto 0);
    hits_o_95 : out std_logic_vector(1 downto 0);
    hits_o_96 : out std_logic_vector(1 downto 0);
    hits_o_97 : out std_logic_vector(1 downto 0);
    hits_o_98 : out std_logic_vector(1 downto 0);
    hits_o_99 : out std_logic_vector(1 downto 0);
    hits_o_100 : out std_logic_vector(1 downto 0);
    hits_o_101 : out std_logic_vector(1 downto 0);
    hits_o_102 : out std_logic_vector(1 downto 0);
    hits_o_103 : out std_logic_vector(1 downto 0);
    hits_o_104 : out std_logic_vector(1 downto 0);
    hits_o_105 : out std_logic_vector(1 downto 0);
    hits_o_106 : out std_logic_vector(1 downto 0);
    hits_o_107 : out std_logic_vector(1 downto 0);
    hits_o_108 : out std_logic_vector(1 downto 0);
    hits_o_109 : out std_logic_vector(1 downto 0);
    hits_o_110 : out std_logic_vector(1 downto 0);
    hits_o_111 : out std_logic_vector(1 downto 0);
    hits_o_112 : out std_logic_vector(1 downto 0);
    hits_o_113 : out std_logic_vector(1 downto 0);
    hits_o_114 : out std_logic_vector(1 downto 0);
    hits_o_115 : out std_logic_vector(1 downto 0);
    hits_o_116 : out std_logic_vector(1 downto 0);
    hits_o_117 : out std_logic_vector(1 downto 0);
    hits_o_118 : out std_logic_vector(1 downto 0);
    hits_o_119 : out std_logic_vector(1 downto 0);
    hits_o_120 : out std_logic_vector(1 downto 0);
    hits_o_121 : out std_logic_vector(1 downto 0);
    hits_o_122 : out std_logic_vector(1 downto 0);
    hits_o_123 : out std_logic_vector(1 downto 0);
    hits_o_124 : out std_logic_vector(1 downto 0);
    hits_o_125 : out std_logic_vector(1 downto 0);
    hits_o_126 : out std_logic_vector(1 downto 0);
    hits_o_127 : out std_logic_vector(1 downto 0);
    hits_o_128 : out std_logic_vector(1 downto 0);
    hits_o_129 : out std_logic_vector(1 downto 0);
    hits_o_130 : out std_logic_vector(1 downto 0);
    hits_o_131 : out std_logic_vector(1 downto 0);
    hits_o_132 : out std_logic_vector(1 downto 0);
    hits_o_133 : out std_logic_vector(1 downto 0);
    hits_o_134 : out std_logic_vector(1 downto 0);
    hits_o_135 : out std_logic_vector(1 downto 0);
    hits_o_136 : out std_logic_vector(1 downto 0);
    hits_o_137 : out std_logic_vector(1 downto 0);
    hits_o_138 : out std_logic_vector(1 downto 0);
    hits_o_139 : out std_logic_vector(1 downto 0);
    hits_o_140 : out std_logic_vector(1 downto 0);
    hits_o_141 : out std_logic_vector(1 downto 0);
    hits_o_142 : out std_logic_vector(1 downto 0);
    hits_o_143 : out std_logic_vector(1 downto 0);
    hits_o_144 : out std_logic_vector(1 downto 0);
    hits_o_145 : out std_logic_vector(1 downto 0);
    hits_o_146 : out std_logic_vector(1 downto 0);
    hits_o_147 : out std_logic_vector(1 downto 0);
    hits_o_148 : out std_logic_vector(1 downto 0);
    hits_o_149 : out std_logic_vector(1 downto 0);
    hits_o_150 : out std_logic_vector(1 downto 0);
    hits_o_151 : out std_logic_vector(1 downto 0);
    hits_o_152 : out std_logic_vector(1 downto 0);
    hits_o_153 : out std_logic_vector(1 downto 0);
    hits_o_154 : out std_logic_vector(1 downto 0);
    hits_o_155 : out std_logic_vector(1 downto 0);
    hits_o_156 : out std_logic_vector(1 downto 0);
    hits_o_157 : out std_logic_vector(1 downto 0);
    hits_o_158 : out std_logic_vector(1 downto 0);
    hits_o_159 : out std_logic_vector(1 downto 0);
    hits_o_160 : out std_logic_vector(1 downto 0);
    hits_o_161 : out std_logic_vector(1 downto 0);
    hits_o_162 : out std_logic_vector(1 downto 0);
    hits_o_163 : out std_logic_vector(1 downto 0);
    hits_o_164 : out std_logic_vector(1 downto 0);
    hits_o_165 : out std_logic_vector(1 downto 0);
    hits_o_166 : out std_logic_vector(1 downto 0);
    hits_o_167 : out std_logic_vector(1 downto 0);
    hits_o_168 : out std_logic_vector(1 downto 0);
    hits_o_169 : out std_logic_vector(1 downto 0);
    hits_o_170 : out std_logic_vector(1 downto 0);
    hits_o_171 : out std_logic_vector(1 downto 0);
    hits_o_172 : out std_logic_vector(1 downto 0);
    hits_o_173 : out std_logic_vector(1 downto 0);
    hits_o_174 : out std_logic_vector(1 downto 0);
    hits_o_175 : out std_logic_vector(1 downto 0);
    hits_o_176 : out std_logic_vector(1 downto 0);
    hits_o_177 : out std_logic_vector(1 downto 0);
    hits_o_178 : out std_logic_vector(1 downto 0);
    hits_o_179 : out std_logic_vector(1 downto 0);
    hits_o_180 : out std_logic_vector(1 downto 0);
    hits_o_181 : out std_logic_vector(1 downto 0);
    hits_o_182 : out std_logic_vector(1 downto 0);
    hits_o_183 : out std_logic_vector(1 downto 0);
    hits_o_184 : out std_logic_vector(1 downto 0);
    hits_o_185 : out std_logic_vector(1 downto 0);
    hits_o_186 : out std_logic_vector(1 downto 0);
    hits_o_187 : out std_logic_vector(1 downto 0);
    hits_o_188 : out std_logic_vector(1 downto 0);
    hits_o_189 : out std_logic_vector(1 downto 0);
    hits_o_190 : out std_logic_vector(1 downto 0);
    hits_o_191 : out std_logic_vector(1 downto 0);
    hits_o_192 : out std_logic_vector(1 downto 0);
    hits_o_193 : out std_logic_vector(1 downto 0);
    hits_o_194 : out std_logic_vector(1 downto 0);
    hits_o_195 : out std_logic_vector(1 downto 0);
    hits_o_196 : out std_logic_vector(1 downto 0);
    hits_o_197 : out std_logic_vector(1 downto 0);
    hits_o_198 : out std_logic_vector(1 downto 0);
    hits_o_199 : out std_logic_vector(1 downto 0);

    -- trigger parameters
    gaps_trigger_en  : in std_logic;
    require_beta     : in std_logic;
    inner_tof_thresh : in std_logic_vector (7 downto 0);
    outer_tof_thresh : in std_logic_vector (7 downto 0);
    total_tof_thresh : in std_logic_vector (7 downto 0);

    busy_i      : in std_logic;
    rb_busy_i   : in std_logic_vector(NUM_RBS-1 downto 0);
    rb_window_i : in std_logic_vector(4 downto 0);

    force_trigger_i : in std_logic;

    trig_sources_o   : out std_logic_vector(15 downto 0);
    pre_trigger_o    : out std_logic;
    global_trigger_o : out std_logic;
    lost_trigger_o   : out std_logic;
    rb_trigger_o     : out std_logic;
    rb_ch_bitmap_o   : out std_logic_vector (NUM_RBS*8-1 downto 0);
    event_cnt_o      : out std_logic_vector (31 downto 0)
    );
end trigger_top;

architecture behavioral of trigger_top is
  signal hits_i : threshold_array_t;
  signal hits_o : threshold_array_t;
begin

  hits_i(0) <= hits_i_0;
  hits_i(1) <= hits_i_1;
  hits_i(2) <= hits_i_2;
  hits_i(3) <= hits_i_3;
  hits_i(4) <= hits_i_4;
  hits_i(5) <= hits_i_5;
  hits_i(6) <= hits_i_6;
  hits_i(7) <= hits_i_7;
  hits_i(8) <= hits_i_8;
  hits_i(9) <= hits_i_9;
  hits_i(10) <= hits_i_10;
  hits_i(11) <= hits_i_11;
  hits_i(12) <= hits_i_12;
  hits_i(13) <= hits_i_13;
  hits_i(14) <= hits_i_14;
  hits_i(15) <= hits_i_15;
  hits_i(16) <= hits_i_16;
  hits_i(17) <= hits_i_17;
  hits_i(18) <= hits_i_18;
  hits_i(19) <= hits_i_19;
  hits_i(20) <= hits_i_20;
  hits_i(21) <= hits_i_21;
  hits_i(22) <= hits_i_22;
  hits_i(23) <= hits_i_23;
  hits_i(24) <= hits_i_24;
  hits_i(25) <= hits_i_25;
  hits_i(26) <= hits_i_26;
  hits_i(27) <= hits_i_27;
  hits_i(28) <= hits_i_28;
  hits_i(29) <= hits_i_29;
  hits_i(30) <= hits_i_30;
  hits_i(31) <= hits_i_31;
  hits_i(32) <= hits_i_32;
  hits_i(33) <= hits_i_33;
  hits_i(34) <= hits_i_34;
  hits_i(35) <= hits_i_35;
  hits_i(36) <= hits_i_36;
  hits_i(37) <= hits_i_37;
  hits_i(38) <= hits_i_38;
  hits_i(39) <= hits_i_39;
  hits_i(40) <= hits_i_40;
  hits_i(41) <= hits_i_41;
  hits_i(42) <= hits_i_42;
  hits_i(43) <= hits_i_43;
  hits_i(44) <= hits_i_44;
  hits_i(45) <= hits_i_45;
  hits_i(46) <= hits_i_46;
  hits_i(47) <= hits_i_47;
  hits_i(48) <= hits_i_48;
  hits_i(49) <= hits_i_49;
  hits_i(50) <= hits_i_50;
  hits_i(51) <= hits_i_51;
  hits_i(52) <= hits_i_52;
  hits_i(53) <= hits_i_53;
  hits_i(54) <= hits_i_54;
  hits_i(55) <= hits_i_55;
  hits_i(56) <= hits_i_56;
  hits_i(57) <= hits_i_57;
  hits_i(58) <= hits_i_58;
  hits_i(59) <= hits_i_59;
  hits_i(60) <= hits_i_60;
  hits_i(61) <= hits_i_61;
  hits_i(62) <= hits_i_62;
  hits_i(63) <= hits_i_63;
  hits_i(64) <= hits_i_64;
  hits_i(65) <= hits_i_65;
  hits_i(66) <= hits_i_66;
  hits_i(67) <= hits_i_67;
  hits_i(68) <= hits_i_68;
  hits_i(69) <= hits_i_69;
  hits_i(70) <= hits_i_70;
  hits_i(71) <= hits_i_71;
  hits_i(72) <= hits_i_72;
  hits_i(73) <= hits_i_73;
  hits_i(74) <= hits_i_74;
  hits_i(75) <= hits_i_75;
  hits_i(76) <= hits_i_76;
  hits_i(77) <= hits_i_77;
  hits_i(78) <= hits_i_78;
  hits_i(79) <= hits_i_79;
  hits_i(80) <= hits_i_80;
  hits_i(81) <= hits_i_81;
  hits_i(82) <= hits_i_82;
  hits_i(83) <= hits_i_83;
  hits_i(84) <= hits_i_84;
  hits_i(85) <= hits_i_85;
  hits_i(86) <= hits_i_86;
  hits_i(87) <= hits_i_87;
  hits_i(88) <= hits_i_88;
  hits_i(89) <= hits_i_89;
  hits_i(90) <= hits_i_90;
  hits_i(91) <= hits_i_91;
  hits_i(92) <= hits_i_92;
  hits_i(93) <= hits_i_93;
  hits_i(94) <= hits_i_94;
  hits_i(95) <= hits_i_95;
  hits_i(96) <= hits_i_96;
  hits_i(97) <= hits_i_97;
  hits_i(98) <= hits_i_98;
  hits_i(99) <= hits_i_99;
  hits_i(100) <= hits_i_100;
  hits_i(101) <= hits_i_101;
  hits_i(102) <= hits_i_102;
  hits_i(103) <= hits_i_103;
  hits_i(104) <= hits_i_104;
  hits_i(105) <= hits_i_105;
  hits_i(106) <= hits_i_106;
  hits_i(107) <= hits_i_107;
  hits_i(108) <= hits_i_108;
  hits_i(109) <= hits_i_109;
  hits_i(110) <= hits_i_110;
  hits_i(111) <= hits_i_111;
  hits_i(112) <= hits_i_112;
  hits_i(113) <= hits_i_113;
  hits_i(114) <= hits_i_114;
  hits_i(115) <= hits_i_115;
  hits_i(116) <= hits_i_116;
  hits_i(117) <= hits_i_117;
  hits_i(118) <= hits_i_118;
  hits_i(119) <= hits_i_119;
  hits_i(120) <= hits_i_120;
  hits_i(121) <= hits_i_121;
  hits_i(122) <= hits_i_122;
  hits_i(123) <= hits_i_123;
  hits_i(124) <= hits_i_124;
  hits_i(125) <= hits_i_125;
  hits_i(126) <= hits_i_126;
  hits_i(127) <= hits_i_127;
  hits_i(128) <= hits_i_128;
  hits_i(129) <= hits_i_129;
  hits_i(130) <= hits_i_130;
  hits_i(131) <= hits_i_131;
  hits_i(132) <= hits_i_132;
  hits_i(133) <= hits_i_133;
  hits_i(134) <= hits_i_134;
  hits_i(135) <= hits_i_135;
  hits_i(136) <= hits_i_136;
  hits_i(137) <= hits_i_137;
  hits_i(138) <= hits_i_138;
  hits_i(139) <= hits_i_139;
  hits_i(140) <= hits_i_140;
  hits_i(141) <= hits_i_141;
  hits_i(142) <= hits_i_142;
  hits_i(143) <= hits_i_143;
  hits_i(144) <= hits_i_144;
  hits_i(145) <= hits_i_145;
  hits_i(146) <= hits_i_146;
  hits_i(147) <= hits_i_147;
  hits_i(148) <= hits_i_148;
  hits_i(149) <= hits_i_149;
  hits_i(150) <= hits_i_150;
  hits_i(151) <= hits_i_151;
  hits_i(152) <= hits_i_152;
  hits_i(153) <= hits_i_153;
  hits_i(154) <= hits_i_154;
  hits_i(155) <= hits_i_155;
  hits_i(156) <= hits_i_156;
  hits_i(157) <= hits_i_157;
  hits_i(158) <= hits_i_158;
  hits_i(159) <= hits_i_159;
  hits_i(160) <= hits_i_160;
  hits_i(161) <= hits_i_161;
  hits_i(162) <= hits_i_162;
  hits_i(163) <= hits_i_163;
  hits_i(164) <= hits_i_164;
  hits_i(165) <= hits_i_165;
  hits_i(166) <= hits_i_166;
  hits_i(167) <= hits_i_167;
  hits_i(168) <= hits_i_168;
  hits_i(169) <= hits_i_169;
  hits_i(170) <= hits_i_170;
  hits_i(171) <= hits_i_171;
  hits_i(172) <= hits_i_172;
  hits_i(173) <= hits_i_173;
  hits_i(174) <= hits_i_174;
  hits_i(175) <= hits_i_175;
  hits_i(176) <= hits_i_176;
  hits_i(177) <= hits_i_177;
  hits_i(178) <= hits_i_178;
  hits_i(179) <= hits_i_179;
  hits_i(180) <= hits_i_180;
  hits_i(181) <= hits_i_181;
  hits_i(182) <= hits_i_182;
  hits_i(183) <= hits_i_183;
  hits_i(184) <= hits_i_184;
  hits_i(185) <= hits_i_185;
  hits_i(186) <= hits_i_186;
  hits_i(187) <= hits_i_187;
  hits_i(188) <= hits_i_188;
  hits_i(189) <= hits_i_189;
  hits_i(190) <= hits_i_190;
  hits_i(191) <= hits_i_191;
  hits_i(192) <= hits_i_192;
  hits_i(193) <= hits_i_193;
  hits_i(194) <= hits_i_194;
  hits_i(195) <= hits_i_195;
  hits_i(196) <= hits_i_196;
  hits_i(197) <= hits_i_197;
  hits_i(198) <= hits_i_198;
  hits_i(199) <= hits_i_199;

  hits_o_0 <= hits_o(0);
  hits_o_1 <= hits_o(1);
  hits_o_2 <= hits_o(2);
  hits_o_3 <= hits_o(3);
  hits_o_4 <= hits_o(4);
  hits_o_5 <= hits_o(5);
  hits_o_6 <= hits_o(6);
  hits_o_7 <= hits_o(7);
  hits_o_8 <= hits_o(8);
  hits_o_9 <= hits_o(9);
  hits_o_10 <= hits_o(10);
  hits_o_11 <= hits_o(11);
  hits_o_12 <= hits_o(12);
  hits_o_13 <= hits_o(13);
  hits_o_14 <= hits_o(14);
  hits_o_15 <= hits_o(15);
  hits_o_16 <= hits_o(16);
  hits_o_17 <= hits_o(17);
  hits_o_18 <= hits_o(18);
  hits_o_19 <= hits_o(19);
  hits_o_20 <= hits_o(20);
  hits_o_21 <= hits_o(21);
  hits_o_22 <= hits_o(22);
  hits_o_23 <= hits_o(23);
  hits_o_24 <= hits_o(24);
  hits_o_25 <= hits_o(25);
  hits_o_26 <= hits_o(26);
  hits_o_27 <= hits_o(27);
  hits_o_28 <= hits_o(28);
  hits_o_29 <= hits_o(29);
  hits_o_30 <= hits_o(30);
  hits_o_31 <= hits_o(31);
  hits_o_32 <= hits_o(32);
  hits_o_33 <= hits_o(33);
  hits_o_34 <= hits_o(34);
  hits_o_35 <= hits_o(35);
  hits_o_36 <= hits_o(36);
  hits_o_37 <= hits_o(37);
  hits_o_38 <= hits_o(38);
  hits_o_39 <= hits_o(39);
  hits_o_40 <= hits_o(40);
  hits_o_41 <= hits_o(41);
  hits_o_42 <= hits_o(42);
  hits_o_43 <= hits_o(43);
  hits_o_44 <= hits_o(44);
  hits_o_45 <= hits_o(45);
  hits_o_46 <= hits_o(46);
  hits_o_47 <= hits_o(47);
  hits_o_48 <= hits_o(48);
  hits_o_49 <= hits_o(49);
  hits_o_50 <= hits_o(50);
  hits_o_51 <= hits_o(51);
  hits_o_52 <= hits_o(52);
  hits_o_53 <= hits_o(53);
  hits_o_54 <= hits_o(54);
  hits_o_55 <= hits_o(55);
  hits_o_56 <= hits_o(56);
  hits_o_57 <= hits_o(57);
  hits_o_58 <= hits_o(58);
  hits_o_59 <= hits_o(59);
  hits_o_60 <= hits_o(60);
  hits_o_61 <= hits_o(61);
  hits_o_62 <= hits_o(62);
  hits_o_63 <= hits_o(63);
  hits_o_64 <= hits_o(64);
  hits_o_65 <= hits_o(65);
  hits_o_66 <= hits_o(66);
  hits_o_67 <= hits_o(67);
  hits_o_68 <= hits_o(68);
  hits_o_69 <= hits_o(69);
  hits_o_70 <= hits_o(70);
  hits_o_71 <= hits_o(71);
  hits_o_72 <= hits_o(72);
  hits_o_73 <= hits_o(73);
  hits_o_74 <= hits_o(74);
  hits_o_75 <= hits_o(75);
  hits_o_76 <= hits_o(76);
  hits_o_77 <= hits_o(77);
  hits_o_78 <= hits_o(78);
  hits_o_79 <= hits_o(79);
  hits_o_80 <= hits_o(80);
  hits_o_81 <= hits_o(81);
  hits_o_82 <= hits_o(82);
  hits_o_83 <= hits_o(83);
  hits_o_84 <= hits_o(84);
  hits_o_85 <= hits_o(85);
  hits_o_86 <= hits_o(86);
  hits_o_87 <= hits_o(87);
  hits_o_88 <= hits_o(88);
  hits_o_89 <= hits_o(89);
  hits_o_90 <= hits_o(90);
  hits_o_91 <= hits_o(91);
  hits_o_92 <= hits_o(92);
  hits_o_93 <= hits_o(93);
  hits_o_94 <= hits_o(94);
  hits_o_95 <= hits_o(95);
  hits_o_96 <= hits_o(96);
  hits_o_97 <= hits_o(97);
  hits_o_98 <= hits_o(98);
  hits_o_99 <= hits_o(99);
  hits_o_100 <= hits_o(100);
  hits_o_101 <= hits_o(101);
  hits_o_102 <= hits_o(102);
  hits_o_103 <= hits_o(103);
  hits_o_104 <= hits_o(104);
  hits_o_105 <= hits_o(105);
  hits_o_106 <= hits_o(106);
  hits_o_107 <= hits_o(107);
  hits_o_108 <= hits_o(108);
  hits_o_109 <= hits_o(109);
  hits_o_110 <= hits_o(110);
  hits_o_111 <= hits_o(111);
  hits_o_112 <= hits_o(112);
  hits_o_113 <= hits_o(113);
  hits_o_114 <= hits_o(114);
  hits_o_115 <= hits_o(115);
  hits_o_116 <= hits_o(116);
  hits_o_117 <= hits_o(117);
  hits_o_118 <= hits_o(118);
  hits_o_119 <= hits_o(119);
  hits_o_120 <= hits_o(120);
  hits_o_121 <= hits_o(121);
  hits_o_122 <= hits_o(122);
  hits_o_123 <= hits_o(123);
  hits_o_124 <= hits_o(124);
  hits_o_125 <= hits_o(125);
  hits_o_126 <= hits_o(126);
  hits_o_127 <= hits_o(127);
  hits_o_128 <= hits_o(128);
  hits_o_129 <= hits_o(129);
  hits_o_130 <= hits_o(130);
  hits_o_131 <= hits_o(131);
  hits_o_132 <= hits_o(132);
  hits_o_133 <= hits_o(133);
  hits_o_134 <= hits_o(134);
  hits_o_135 <= hits_o(135);
  hits_o_136 <= hits_o(136);
  hits_o_137 <= hits_o(137);
  hits_o_138 <= hits_o(138);
  hits_o_139 <= hits_o(139);
  hits_o_140 <= hits_o(140);
  hits_o_141 <= hits_o(141);
  hits_o_142 <= hits_o(142);
  hits_o_143 <= hits_o(143);
  hits_o_144 <= hits_o(144);
  hits_o_145 <= hits_o(145);
  hits_o_146 <= hits_o(146);
  hits_o_147 <= hits_o(147);
  hits_o_148 <= hits_o(148);
  hits_o_149 <= hits_o(149);
  hits_o_150 <= hits_o(150);
  hits_o_151 <= hits_o(151);
  hits_o_152 <= hits_o(152);
  hits_o_153 <= hits_o(153);
  hits_o_154 <= hits_o(154);
  hits_o_155 <= hits_o(155);
  hits_o_156 <= hits_o(156);
  hits_o_157 <= hits_o(157);
  hits_o_158 <= hits_o(158);
  hits_o_159 <= hits_o(159);
  hits_o_160 <= hits_o(160);
  hits_o_161 <= hits_o(161);
  hits_o_162 <= hits_o(162);
  hits_o_163 <= hits_o(163);
  hits_o_164 <= hits_o(164);
  hits_o_165 <= hits_o(165);
  hits_o_166 <= hits_o(166);
  hits_o_167 <= hits_o(167);
  hits_o_168 <= hits_o(168);
  hits_o_169 <= hits_o(169);
  hits_o_170 <= hits_o(170);
  hits_o_171 <= hits_o(171);
  hits_o_172 <= hits_o(172);
  hits_o_173 <= hits_o(173);
  hits_o_174 <= hits_o(174);
  hits_o_175 <= hits_o(175);
  hits_o_176 <= hits_o(176);
  hits_o_177 <= hits_o(177);
  hits_o_178 <= hits_o(178);
  hits_o_179 <= hits_o(179);
  hits_o_180 <= hits_o(180);
  hits_o_181 <= hits_o(181);
  hits_o_182 <= hits_o(182);
  hits_o_183 <= hits_o(183);
  hits_o_184 <= hits_o(184);
  hits_o_185 <= hits_o(185);
  hits_o_186 <= hits_o(186);
  hits_o_187 <= hits_o(187);
  hits_o_188 <= hits_o(188);
  hits_o_189 <= hits_o(189);
  hits_o_190 <= hits_o(190);
  hits_o_191 <= hits_o(191);
  hits_o_192 <= hits_o(192);
  hits_o_193 <= hits_o(193);
  hits_o_194 <= hits_o(194);
  hits_o_195 <= hits_o(195);
  hits_o_196 <= hits_o(196);
  hits_o_197 <= hits_o(197);
  hits_o_198 <= hits_o(198);
  hits_o_199 <= hits_o(199);


  trigger_2: entity work.trigger
    generic map (
      DEBUG => DEBUG)
    port map (
      clk                       => clk,
      reset                     => reset,
      event_cnt_reset           => event_cnt_reset,
      any_hit_trigger_is_global => any_hit_trigger_is_global,
      track_trigger_is_global   => track_trigger_is_global,
      track_central_is_global   => track_central_is_global,
      any_hit_trigger_prescale  => any_hit_trigger_prescale,
      track_trigger_prescale    => track_trigger_prescale,
      track_central_prescale    => track_central_prescale,
      hit_thresh                => hit_thresh,
      read_all_channels         => read_all_channels,
      hits_i                    => hits_i,
      hits_o                    => hits_o,
      gaps_trigger_en           => gaps_trigger_en,
      require_beta              => require_beta,
      inner_tof_thresh          => inner_tof_thresh,
      outer_tof_thresh          => outer_tof_thresh,
      total_tof_thresh          => total_tof_thresh,
      busy_i                    => busy_i,
      rb_busy_i                 => rb_busy_i,
      rb_window_i               => rb_window_i,
      force_trigger_i           => force_trigger_i,
      trig_sources_o            => trig_sources_o,
      pre_trigger_o             => pre_trigger_o,
      global_trigger_o          => global_trigger_o,
      lost_trigger_o            => lost_trigger_o,
      rb_trigger_o              => rb_trigger_o,
      rb_ch_bitmap_o            => rb_ch_bitmap_o,
      event_cnt_o               => event_cnt_o);

end behavioral;
