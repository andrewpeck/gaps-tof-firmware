library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.types_pkg.all;
use work.mt_types.all;
use work.constants.all;
use work.components.all;

entity rb_map is
  port(
    clock          : in  std_logic;
    hits_bitmap_i  : in  channel_bitmask_t := (others => '0');
    rb_ch_bitmap_o : out std_logic_vector (NUM_RBS*8-1 downto 0) -- 399 downto 0
    );
end rb_map;

architecture behavioral of rb_map is
begin

  -- rb_ch_bitmap_o(399 downto 0) <= hits_bitmap_i(199 downto 0);
  --
  -- this file maps from LTB channels on the right hand side, to readout board
  -- channels on the left hand side.
  --
  -- so e.g. LTB input 0 (DSI1, J1, BIT1) is represented by hits_bitmap_i(0)
  --

  --START: autoinsert mapping

  rb_ch_bitmap_o(196) <= hits_bitmap_i( 61); -- {:station "cube", :ltb-harting 2, :paddle-number 1, :ltb-num+channel {:board 8, :ch 11}, :rb-num+channel {:board 15, :ch 5}, :dsi-slot 2, :panel-number 1, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(196) <= hits_bitmap_i( 60); -- {:station "cube", :ltb-harting 2, :paddle-number 2, :ltb-num+channel {:board 8, :ch 9}, :rb-num+channel {:board 16, :ch 5}, :dsi-slot 2, :panel-number 1, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(194) <= hits_bitmap_i( 59); -- {:station "cube", :ltb-harting 2, :paddle-number 3, :ltb-num+channel {:board 8, :ch 7}, :rb-num+channel {:board 15, :ch 3}, :dsi-slot 2, :panel-number 1, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(194) <= hits_bitmap_i( 58); -- {:station "cube", :ltb-harting 2, :paddle-number 4, :ltb-num+channel {:board 8, :ch 5}, :rb-num+channel {:board 16, :ch 3}, :dsi-slot 2, :panel-number 1, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(192) <= hits_bitmap_i( 57); -- {:station "cube", :ltb-harting 2, :paddle-number 5, :ltb-num+channel {:board 8, :ch 3}, :rb-num+channel {:board 15, :ch 1}, :dsi-slot 2, :panel-number 1, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(192) <= hits_bitmap_i( 56); -- {:station "cube", :ltb-harting 2, :paddle-number 6, :ltb-num+channel {:board 8, :ch 1}, :rb-num+channel {:board 16, :ch 1}, :dsi-slot 2, :panel-number 1, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(327) <= hits_bitmap_i(127); -- {:station "cube", :ltb-harting 0, :paddle-number 7, :ltb-num+channel {:board 16, :ch 16}, :rb-num+channel {:board 32, :ch 8}, :dsi-slot 4, :panel-number 1, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(327) <= hits_bitmap_i(126); -- {:station "cube", :ltb-harting 0, :paddle-number 8, :ltb-num+channel {:board 16, :ch 14}, :rb-num+channel {:board 31, :ch 8}, :dsi-slot 4, :panel-number 1, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(325) <= hits_bitmap_i(125); -- {:station "cube", :ltb-harting 0, :paddle-number 9, :ltb-num+channel {:board 16, :ch 12}, :rb-num+channel {:board 32, :ch 6}, :dsi-slot 4, :panel-number 1, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(325) <= hits_bitmap_i(124); -- {:station "cube", :ltb-harting 0, :paddle-number 10, :ltb-num+channel {:board 16, :ch 10}, :rb-num+channel {:board 31, :ch 6}, :dsi-slot 4, :panel-number 1, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(323) <= hits_bitmap_i(123); -- {:station "cube", :ltb-harting 0, :paddle-number 11, :ltb-num+channel {:board 16, :ch 8}, :rb-num+channel {:board 32, :ch 4}, :dsi-slot 4, :panel-number 1, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(323) <= hits_bitmap_i(122); -- {:station "cube", :ltb-harting 0, :paddle-number 12, :ltb-num+channel {:board 16, :ch 6}, :rb-num+channel {:board 31, :ch 4}, :dsi-slot 4, :panel-number 1, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(225) <= hits_bitmap_i( 72); -- {:station "cube_bot", :ltb-harting 4, :paddle-number 13, :ltb-num+channel {:board 10, :ch 2}, :rb-num+channel {:board 19, :ch 2}, :dsi-slot 2, :panel-number 2, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(225) <= hits_bitmap_i( 73); -- {:station "cube_bot", :ltb-harting 4, :paddle-number 14, :ltb-num+channel {:board 10, :ch 4}, :rb-num+channel {:board 20, :ch 2}, :dsi-slot 2, :panel-number 2, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(227) <= hits_bitmap_i( 74); -- {:station "cube_bot", :ltb-harting 4, :paddle-number 15, :ltb-num+channel {:board 10, :ch 6}, :rb-num+channel {:board 19, :ch 4}, :dsi-slot 2, :panel-number 2, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(227) <= hits_bitmap_i( 75); -- {:station "cube_bot", :ltb-harting 4, :paddle-number 16, :ltb-num+channel {:board 10, :ch 8}, :rb-num+channel {:board 20, :ch 4}, :dsi-slot 2, :panel-number 2, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(229) <= hits_bitmap_i( 76); -- {:station "cube_bot", :ltb-harting 4, :paddle-number 17, :ltb-num+channel {:board 10, :ch 10}, :rb-num+channel {:board 19, :ch 6}, :dsi-slot 2, :panel-number 2, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(229) <= hits_bitmap_i( 77); -- {:station "cube_bot", :ltb-harting 4, :paddle-number 18, :ltb-num+channel {:board 10, :ch 12}, :rb-num+channel {:board 20, :ch 6}, :dsi-slot 2, :panel-number 2, :paddle-end :A, :rb-harting 4, :rat-number 10}
  rb_ch_bitmap_o(290) <= hits_bitmap_i(106); -- {:station "cube_bot", :ltb-harting 3, :paddle-number 19, :ltb-num+channel {:board 14, :ch 5}, :rb-num+channel {:board 28, :ch 3}, :dsi-slot 3, :panel-number 2, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(290) <= hits_bitmap_i(107); -- {:station "cube_bot", :ltb-harting 3, :paddle-number 20, :ltb-num+channel {:board 14, :ch 7}, :rb-num+channel {:board 27, :ch 3}, :dsi-slot 3, :panel-number 2, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(292) <= hits_bitmap_i(108); -- {:station "cube_bot", :ltb-harting 3, :paddle-number 21, :ltb-num+channel {:board 14, :ch 9}, :rb-num+channel {:board 28, :ch 5}, :dsi-slot 3, :panel-number 2, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(292) <= hits_bitmap_i(109); -- {:station "cube_bot", :ltb-harting 3, :paddle-number 22, :ltb-num+channel {:board 14, :ch 11}, :rb-num+channel {:board 27, :ch 5}, :dsi-slot 3, :panel-number 2, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(294) <= hits_bitmap_i(110); -- {:station "cube_bot", :ltb-harting 3, :paddle-number 23, :ltb-num+channel {:board 14, :ch 13}, :rb-num+channel {:board 28, :ch 7}, :dsi-slot 3, :panel-number 2, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(294) <= hits_bitmap_i(111); -- {:station "cube_bot", :ltb-harting 3, :paddle-number 24, :ltb-num+channel {:board 14, :ch 15}, :rb-num+channel {:board 27, :ch 7}, :dsi-slot 3, :panel-number 2, :paddle-end :A, :rb-harting 3, :rat-number 14}
  rb_ch_bitmap_o(199) <= hits_bitmap_i( 62); -- {:station "cube", :ltb-harting 2, :paddle-number 25, :ltb-num+channel {:board 8, :ch 14}, :rb-num+channel {:board 16, :ch 8}, :dsi-slot 2, :panel-number 3, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(199) <= hits_bitmap_i( 63); -- {:station "cube", :ltb-harting 2, :paddle-number 26, :ltb-num+channel {:board 8, :ch 16}, :rb-num+channel {:board 15, :ch 8}, :dsi-slot 2, :panel-number 3, :paddle-end :A, :rb-harting 2, :rat-number 8}
  rb_ch_bitmap_o(213) <= hits_bitmap_i( 69); -- {:station "cube", :ltb-harting 3, :paddle-number 27, :ltb-num+channel {:board 9, :ch 12}, :rb-num+channel {:board 18, :ch 6}, :dsi-slot 2, :panel-number 3, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(213) <= hits_bitmap_i( 68); -- {:station "cube", :ltb-harting 3, :paddle-number 28, :ltb-num+channel {:board 9, :ch 10}, :rb-num+channel {:board 17, :ch 6}, :dsi-slot 2, :panel-number 3, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(211) <= hits_bitmap_i( 67); -- {:station "cube", :ltb-harting 3, :paddle-number 29, :ltb-num+channel {:board 9, :ch 8}, :rb-num+channel {:board 18, :ch 4}, :dsi-slot 2, :panel-number 3, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(211) <= hits_bitmap_i( 66); -- {:station "cube", :ltb-harting 3, :paddle-number 30, :ltb-num+channel {:board 9, :ch 6}, :rb-num+channel {:board 17, :ch 4}, :dsi-slot 2, :panel-number 3, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(209) <= hits_bitmap_i( 65); -- {:station "cube", :ltb-harting 3, :paddle-number 31, :ltb-num+channel {:board 9, :ch 4}, :rb-num+channel {:board 18, :ch 2}, :dsi-slot 2, :panel-number 3, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(209) <= hits_bitmap_i( 64); -- {:station "cube", :ltb-harting 3, :paddle-number 32, :ltb-num+channel {:board 9, :ch 2}, :rb-num+channel {:board 17, :ch 2}, :dsi-slot 2, :panel-number 3, :paddle-end :A, :rb-harting 3, :rat-number 9}
  rb_ch_bitmap_o(263) <= hits_bitmap_i( 92); -- {:station "cube", :ltb-harting 1, :paddle-number 33, :ltb-num+channel {:board 12, :ch 10}, :rb-num+channel {:board 24, :ch 8}, :dsi-slot 3, :panel-number 4, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(263) <= hits_bitmap_i( 91); -- {:station "cube", :ltb-harting 1, :paddle-number 34, :ltb-num+channel {:board 12, :ch 8}, :rb-num+channel {:board 23, :ch 8}, :dsi-slot 3, :panel-number 4, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(261) <= hits_bitmap_i( 93); -- {:station "cube", :ltb-harting 1, :paddle-number 35, :ltb-num+channel {:board 12, :ch 12}, :rb-num+channel {:board 24, :ch 6}, :dsi-slot 3, :panel-number 4, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(261) <= hits_bitmap_i( 90); -- {:station "cube", :ltb-harting 1, :paddle-number 36, :ltb-num+channel {:board 12, :ch 6}, :rb-num+channel {:board 23, :ch 6}, :dsi-slot 3, :panel-number 4, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(259) <= hits_bitmap_i( 94); -- {:station "cube", :ltb-harting 1, :paddle-number 37, :ltb-num+channel {:board 12, :ch 14}, :rb-num+channel {:board 24, :ch 4}, :dsi-slot 3, :panel-number 4, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(259) <= hits_bitmap_i( 89); -- {:station "cube", :ltb-harting 1, :paddle-number 38, :ltb-num+channel {:board 12, :ch 4}, :rb-num+channel {:board 23, :ch 4}, :dsi-slot 3, :panel-number 4, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(257) <= hits_bitmap_i( 95); -- {:station "cube", :ltb-harting 1, :paddle-number 39, :ltb-num+channel {:board 12, :ch 16}, :rb-num+channel {:board 24, :ch 2}, :dsi-slot 3, :panel-number 4, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(257) <= hits_bitmap_i( 88); -- {:station "cube", :ltb-harting 1, :paddle-number 40, :ltb-num+channel {:board 12, :ch 2}, :rb-num+channel {:board 23, :ch 2}, :dsi-slot 3, :panel-number 4, :paddle-end :A, :rb-harting 1, :rat-number 12}
  rb_ch_bitmap_o(321) <= hits_bitmap_i(121); -- {:station "cube", :ltb-harting 0, :paddle-number 41, :ltb-num+channel {:board 16, :ch 4}, :rb-num+channel {:board 32, :ch 2}, :dsi-slot 4, :panel-number 5, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(321) <= hits_bitmap_i(120); -- {:station "cube", :ltb-harting 0, :paddle-number 42, :ltb-num+channel {:board 16, :ch 2}, :rb-num+channel {:board 31, :ch 2}, :dsi-slot 4, :panel-number 5, :paddle-end :A, :rb-harting 0, :rat-number 16}
  rb_ch_bitmap_o(307) <= hits_bitmap_i(114); -- {:station "cube", :ltb-harting 4, :paddle-number 43, :ltb-num+channel {:board 15, :ch 6}, :rb-num+channel {:board 30, :ch 4}, :dsi-slot 3, :panel-number 5, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(307) <= hits_bitmap_i(115); -- {:station "cube", :ltb-harting 4, :paddle-number 44, :ltb-num+channel {:board 15, :ch 8}, :rb-num+channel {:board 29, :ch 4}, :dsi-slot 3, :panel-number 5, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(309) <= hits_bitmap_i(116); -- {:station "cube", :ltb-harting 4, :paddle-number 45, :ltb-num+channel {:board 15, :ch 10}, :rb-num+channel {:board 30, :ch 6}, :dsi-slot 3, :panel-number 5, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(309) <= hits_bitmap_i(117); -- {:station "cube", :ltb-harting 4, :paddle-number 46, :ltb-num+channel {:board 15, :ch 12}, :rb-num+channel {:board 29, :ch 6}, :dsi-slot 3, :panel-number 5, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(311) <= hits_bitmap_i(118); -- {:station "cube", :ltb-harting 4, :paddle-number 47, :ltb-num+channel {:board 15, :ch 14}, :rb-num+channel {:board 30, :ch 8}, :dsi-slot 3, :panel-number 5, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(311) <= hits_bitmap_i(119); -- {:station "cube", :ltb-harting 4, :paddle-number 48, :ltb-num+channel {:board 15, :ch 16}, :rb-num+channel {:board 29, :ch 8}, :dsi-slot 3, :panel-number 5, :paddle-end :A, :rb-harting 4, :rat-number 15}
  rb_ch_bitmap_o(375) <= hits_bitmap_i(148); -- {:station "cube", :ltb-harting 3, :paddle-number 49, :ltb-num+channel {:board 19, :ch 10}, :rb-num+channel {:board 38, :ch 8}, :dsi-slot 4, :panel-number 6, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(375) <= hits_bitmap_i(147); -- {:station "cube", :ltb-harting 3, :paddle-number 50, :ltb-num+channel {:board 19, :ch 8}, :rb-num+channel {:board 37, :ch 8}, :dsi-slot 4, :panel-number 6, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(373) <= hits_bitmap_i(149); -- {:station "cube", :ltb-harting 3, :paddle-number 51, :ltb-num+channel {:board 19, :ch 12}, :rb-num+channel {:board 38, :ch 6}, :dsi-slot 4, :panel-number 6, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(373) <= hits_bitmap_i(146); -- {:station "cube", :ltb-harting 3, :paddle-number 52, :ltb-num+channel {:board 19, :ch 6}, :rb-num+channel {:board 37, :ch 6}, :dsi-slot 4, :panel-number 6, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(371) <= hits_bitmap_i(150); -- {:station "cube", :ltb-harting 3, :paddle-number 53, :ltb-num+channel {:board 19, :ch 14}, :rb-num+channel {:board 38, :ch 4}, :dsi-slot 4, :panel-number 6, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(371) <= hits_bitmap_i(145); -- {:station "cube", :ltb-harting 3, :paddle-number 54, :ltb-num+channel {:board 19, :ch 4}, :rb-num+channel {:board 37, :ch 4}, :dsi-slot 4, :panel-number 6, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(369) <= hits_bitmap_i(151); -- {:station "cube", :ltb-harting 3, :paddle-number 55, :ltb-num+channel {:board 19, :ch 16}, :rb-num+channel {:board 38, :ch 2}, :dsi-slot 4, :panel-number 6, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(369) <= hits_bitmap_i(144); -- {:station "cube", :ltb-harting 3, :paddle-number 56, :ltb-num+channel {:board 19, :ch 2}, :rb-num+channel {:board 37, :ch 2}, :dsi-slot 4, :panel-number 6, :paddle-end :A, :rb-harting 3, :rat-number 19}
  rb_ch_bitmap_o(241) <= hits_bitmap_i( 81); -- {:station "cube_corner", :ltb-harting 0, :paddle-number 57, :ltb-num+channel {:board 11, :ch 4}, :rb-num+channel {:board 21, :ch 2}, :dsi-slot 3, :panel-number "E-X045", :paddle-end :A, :rb-harting 0, :rat-number 11}
  rb_ch_bitmap_o(279) <= hits_bitmap_i(102); -- {:station "cube_corner", :ltb-harting 2, :paddle-number 58, :ltb-num+channel {:board 13, :ch 14}, :rb-num+channel {:board 25, :ch 8}, :dsi-slot 3, :panel-number "E-X135", :paddle-end :A, :rb-harting 2, :rat-number 13}
  rb_ch_bitmap_o(337) <= hits_bitmap_i(129); -- {:station "cube_corner", :ltb-harting 1, :paddle-number 59, :ltb-num+channel {:board 17, :ch 4}, :rb-num+channel {:board 33, :ch 2}, :dsi-slot 4, :panel-number "E-X225", :paddle-end :A, :rb-harting 1, :rat-number 17}
  rb_ch_bitmap_o(183) <= hits_bitmap_i( 54); -- {:station "cube_corner", :ltb-harting 1, :paddle-number 60, :ltb-num+channel {:board 7, :ch 14}, :rb-num+channel {:board 13, :ch 8}, :dsi-slot 2, :panel-number "E-X315", :paddle-end :A, :rb-harting 1, :rat-number 7}
  rb_ch_bitmap_o( 84) <= hits_bitmap_i(  5); -- {:station "umbrella", :ltb-harting 0, :paddle-number 61, :ltb-num+channel {:board 1, :ch 11}, :rb-num+channel {:board 2, :ch 5}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 84) <= hits_bitmap_i(  4); -- {:station "umbrella", :ltb-harting 0, :paddle-number 62, :ltb-num+channel {:board 1, :ch 9}, :rb-num+channel {:board 1, :ch 5}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 82) <= hits_bitmap_i(  3); -- {:station "umbrella", :ltb-harting 0, :paddle-number 63, :ltb-num+channel {:board 1, :ch 7}, :rb-num+channel {:board 2, :ch 3}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 82) <= hits_bitmap_i(  2); -- {:station "umbrella", :ltb-harting 0, :paddle-number 64, :ltb-num+channel {:board 1, :ch 5}, :rb-num+channel {:board 1, :ch 3}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 80) <= hits_bitmap_i(  1); -- {:station "umbrella", :ltb-harting 0, :paddle-number 65, :ltb-num+channel {:board 1, :ch 3}, :rb-num+channel {:board 2, :ch 1}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 80) <= hits_bitmap_i(  0); -- {:station "umbrella", :ltb-harting 0, :paddle-number 66, :ltb-num+channel {:board 1, :ch 1}, :rb-num+channel {:board 1, :ch 1}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 97) <= hits_bitmap_i(  8); -- {:station "umbrella", :ltb-harting 1, :paddle-number 67, :ltb-num+channel {:board 2, :ch 2}, :rb-num+channel {:board 3, :ch 2}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 97) <= hits_bitmap_i(  9); -- {:station "umbrella", :ltb-harting 1, :paddle-number 68, :ltb-num+channel {:board 2, :ch 4}, :rb-num+channel {:board 4, :ch 2}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 99) <= hits_bitmap_i( 10); -- {:station "umbrella", :ltb-harting 1, :paddle-number 69, :ltb-num+channel {:board 2, :ch 6}, :rb-num+channel {:board 3, :ch 4}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 99) <= hits_bitmap_i( 11); -- {:station "umbrella", :ltb-harting 1, :paddle-number 70, :ltb-num+channel {:board 2, :ch 8}, :rb-num+channel {:board 4, :ch 4}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o(101) <= hits_bitmap_i( 12); -- {:station "umbrella", :ltb-harting 1, :paddle-number 71, :ltb-num+channel {:board 2, :ch 10}, :rb-num+channel {:board 3, :ch 6}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o(101) <= hits_bitmap_i( 13); -- {:station "umbrella", :ltb-harting 1, :paddle-number 72, :ltb-num+channel {:board 2, :ch 12}, :rb-num+channel {:board 4, :ch 6}, :dsi-slot 1, :panel-number 7, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o( 86) <= hits_bitmap_i(  6); -- {:station "umbrella", :ltb-harting 0, :paddle-number 73, :ltb-num+channel {:board 1, :ch 13}, :rb-num+channel {:board 2, :ch 7}, :dsi-slot 1, :panel-number 8, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o( 86) <= hits_bitmap_i(  7); -- {:station "umbrella", :ltb-harting 0, :paddle-number 74, :ltb-num+channel {:board 1, :ch 15}, :rb-num+channel {:board 1, :ch 7}, :dsi-slot 1, :panel-number 8, :paddle-end :A, :rb-harting 0, :rat-number 1}
  rb_ch_bitmap_o(112) <= hits_bitmap_i( 16); -- {:station "umbrella", :ltb-harting 2, :paddle-number 75, :ltb-num+channel {:board 3, :ch 1}, :rb-num+channel {:board 5, :ch 1}, :dsi-slot 1, :panel-number 8, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o(112) <= hits_bitmap_i( 17); -- {:station "umbrella", :ltb-harting 2, :paddle-number 76, :ltb-num+channel {:board 3, :ch 3}, :rb-num+channel {:board 6, :ch 1}, :dsi-slot 1, :panel-number 8, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o(114) <= hits_bitmap_i( 18); -- {:station "umbrella", :ltb-harting 2, :paddle-number 77, :ltb-num+channel {:board 3, :ch 5}, :rb-num+channel {:board 5, :ch 3}, :dsi-slot 1, :panel-number 8, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o(114) <= hits_bitmap_i( 19); -- {:station "umbrella", :ltb-harting 2, :paddle-number 78, :ltb-num+channel {:board 3, :ch 7}, :rb-num+channel {:board 6, :ch 3}, :dsi-slot 1, :panel-number 8, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o(150) <= hits_bitmap_i( 39); -- {:station "umbrella", :ltb-harting 4, :paddle-number 79, :ltb-num+channel {:board 5, :ch 15}, :rb-num+channel {:board 9, :ch 7}, :dsi-slot 1, :panel-number 9, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o(150) <= hits_bitmap_i( 38); -- {:station "umbrella", :ltb-harting 4, :paddle-number 80, :ltb-num+channel {:board 5, :ch 13}, :rb-num+channel {:board 10, :ch 7}, :dsi-slot 1, :panel-number 9, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o(148) <= hits_bitmap_i( 37); -- {:station "umbrella", :ltb-harting 4, :paddle-number 81, :ltb-num+channel {:board 5, :ch 11}, :rb-num+channel {:board 9, :ch 5}, :dsi-slot 1, :panel-number 9, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o(148) <= hits_bitmap_i( 36); -- {:station "umbrella", :ltb-harting 4, :paddle-number 82, :ltb-num+channel {:board 5, :ch 9}, :rb-num+channel {:board 10, :ch 5}, :dsi-slot 1, :panel-number 9, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o(146) <= hits_bitmap_i( 35); -- {:station "umbrella", :ltb-harting 4, :paddle-number 83, :ltb-num+channel {:board 5, :ch 7}, :rb-num+channel {:board 9, :ch 3}, :dsi-slot 1, :panel-number 9, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o(146) <= hits_bitmap_i( 34); -- {:station "umbrella", :ltb-harting 4, :paddle-number 84, :ltb-num+channel {:board 5, :ch 5}, :rb-num+channel {:board 10, :ch 3}, :dsi-slot 1, :panel-number 9, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o(144) <= hits_bitmap_i( 33); -- {:station "umbrella", :ltb-harting 4, :paddle-number 85, :ltb-num+channel {:board 5, :ch 3}, :rb-num+channel {:board 10, :ch 1}, :dsi-slot 1, :panel-number 10, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o(144) <= hits_bitmap_i( 32); -- {:station "umbrella", :ltb-harting 4, :paddle-number 86, :ltb-num+channel {:board 5, :ch 1}, :rb-num+channel {:board 9, :ch 1}, :dsi-slot 1, :panel-number 10, :paddle-end :A, :rb-harting 4, :rat-number 5}
  rb_ch_bitmap_o(134) <= hits_bitmap_i( 31); -- {:station "umbrella", :ltb-harting 3, :paddle-number 87, :ltb-num+channel {:board 4, :ch 15}, :rb-num+channel {:board 7, :ch 7}, :dsi-slot 1, :panel-number 10, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o(134) <= hits_bitmap_i( 30); -- {:station "umbrella", :ltb-harting 3, :paddle-number 88, :ltb-num+channel {:board 4, :ch 13}, :rb-num+channel {:board 8, :ch 7}, :dsi-slot 1, :panel-number 10, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o(132) <= hits_bitmap_i( 29); -- {:station "umbrella", :ltb-harting 3, :paddle-number 89, :ltb-num+channel {:board 4, :ch 11}, :rb-num+channel {:board 7, :ch 5}, :dsi-slot 1, :panel-number 10, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o(132) <= hits_bitmap_i( 28); -- {:station "umbrella", :ltb-harting 3, :paddle-number 90, :ltb-num+channel {:board 4, :ch 9}, :rb-num+channel {:board 8, :ch 5}, :dsi-slot 1, :panel-number 10, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o(103) <= hits_bitmap_i( 14); -- {:station "umbrella", :ltb-harting 1, :paddle-number 91, :ltb-num+channel {:board 2, :ch 14}, :rb-num+channel {:board 4, :ch 8}, :dsi-slot 1, :panel-number 11, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o(103) <= hits_bitmap_i( 15); -- {:station "umbrella", :ltb-harting 1, :paddle-number 92, :ltb-num+channel {:board 2, :ch 16}, :rb-num+channel {:board 3, :ch 8}, :dsi-slot 1, :panel-number 11, :paddle-end :A, :rb-harting 1, :rat-number 2}
  rb_ch_bitmap_o(128) <= hits_bitmap_i( 24); -- {:station "umbrella", :ltb-harting 3, :paddle-number 93, :ltb-num+channel {:board 4, :ch 1}, :rb-num+channel {:board 7, :ch 1}, :dsi-slot 1, :panel-number 11, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o(128) <= hits_bitmap_i( 25); -- {:station "umbrella", :ltb-harting 3, :paddle-number 94, :ltb-num+channel {:board 4, :ch 3}, :rb-num+channel {:board 8, :ch 1}, :dsi-slot 1, :panel-number 11, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o(130) <= hits_bitmap_i( 26); -- {:station "umbrella", :ltb-harting 3, :paddle-number 95, :ltb-num+channel {:board 4, :ch 5}, :rb-num+channel {:board 7, :ch 3}, :dsi-slot 1, :panel-number 11, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o(130) <= hits_bitmap_i( 27); -- {:station "umbrella", :ltb-harting 3, :paddle-number 96, :ltb-num+channel {:board 4, :ch 7}, :rb-num+channel {:board 8, :ch 3}, :dsi-slot 1, :panel-number 11, :paddle-end :A, :rb-harting 3, :rat-number 4}
  rb_ch_bitmap_o(166) <= hits_bitmap_i( 47); -- {:station "umbrella", :ltb-harting 0, :paddle-number 97, :ltb-num+channel {:board 6, :ch 15}, :rb-num+channel {:board 11, :ch 7}, :dsi-slot 2, :panel-number 12, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o(166) <= hits_bitmap_i( 46); -- {:station "umbrella", :ltb-harting 0, :paddle-number 98, :ltb-num+channel {:board 6, :ch 13}, :rb-num+channel {:board 12, :ch 7}, :dsi-slot 2, :panel-number 12, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o(164) <= hits_bitmap_i( 45); -- {:station "umbrella", :ltb-harting 0, :paddle-number 99, :ltb-num+channel {:board 6, :ch 11}, :rb-num+channel {:board 11, :ch 5}, :dsi-slot 2, :panel-number 12, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o(164) <= hits_bitmap_i( 44); -- {:station "umbrella", :ltb-harting 0, :paddle-number 100, :ltb-num+channel {:board 6, :ch 9}, :rb-num+channel {:board 12, :ch 5}, :dsi-slot 2, :panel-number 12, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o(162) <= hits_bitmap_i( 43); -- {:station "umbrella", :ltb-harting 0, :paddle-number 101, :ltb-num+channel {:board 6, :ch 7}, :rb-num+channel {:board 11, :ch 3}, :dsi-slot 2, :panel-number 12, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o(162) <= hits_bitmap_i( 42); -- {:station "umbrella", :ltb-harting 0, :paddle-number 102, :ltb-num+channel {:board 6, :ch 5}, :rb-num+channel {:board 12, :ch 3}, :dsi-slot 2, :panel-number 12, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o(160) <= hits_bitmap_i( 41); -- {:station "umbrella", :ltb-harting 0, :paddle-number 103, :ltb-num+channel {:board 6, :ch 3}, :rb-num+channel {:board 12, :ch 1}, :dsi-slot 2, :panel-number 13, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o(160) <= hits_bitmap_i( 40); -- {:station "umbrella", :ltb-harting 0, :paddle-number 104, :ltb-num+channel {:board 6, :ch 1}, :rb-num+channel {:board 11, :ch 1}, :dsi-slot 2, :panel-number 13, :paddle-end :A, :rb-harting 0, :rat-number 6}
  rb_ch_bitmap_o(118) <= hits_bitmap_i( 23); -- {:station "umbrella", :ltb-harting 2, :paddle-number 105, :ltb-num+channel {:board 3, :ch 15}, :rb-num+channel {:board 5, :ch 7}, :dsi-slot 1, :panel-number 13, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o(118) <= hits_bitmap_i( 22); -- {:station "umbrella", :ltb-harting 2, :paddle-number 106, :ltb-num+channel {:board 3, :ch 13}, :rb-num+channel {:board 6, :ch 7}, :dsi-slot 1, :panel-number 13, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o(116) <= hits_bitmap_i( 21); -- {:station "umbrella", :ltb-harting 2, :paddle-number 107, :ltb-num+channel {:board 3, :ch 11}, :rb-num+channel {:board 5, :ch 5}, :dsi-slot 1, :panel-number 13, :paddle-end :A, :rb-harting 2, :rat-number 3}
  rb_ch_bitmap_o(116) <= hits_bitmap_i( 20); -- {:station "umbrella", :ltb-harting 2, :paddle-number 108, :ltb-num+channel {:board 3, :ch 9}, :rb-num+channel {:board 6, :ch 5}, :dsi-slot 1, :panel-number 13, :paddle-end :A, :rb-harting 2, :rat-number 3}
-- Failed to map                             -- {:station "cortina", :ltb-harting 3, :paddle-number 109, :ltb-num+channel {:board 9, :ch 16}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 14, :paddle-end :A, :rb-harting 3, :rat-number 9}
-- Failed to map                             -- {:station "cortina", :ltb-harting 3, :paddle-number 110, :ltb-num+channel {:board 9, :ch 14}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 14, :paddle-end :A, :rb-harting 3, :rat-number 9}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 111, :ltb-num+channel {:board 10, :ch 16}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 14, :paddle-end :A, :rb-harting 4, :rat-number 10}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 112, :ltb-num+channel {:board 10, :ch 14}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 14, :paddle-end :A, :rb-harting 4, :rat-number 10}
-- Failed to map                             -- {:station "cortina", :ltb-harting 0, :paddle-number 113, :ltb-num+channel {:board 11, :ch 10}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 14, :paddle-end :A, :rb-harting 0, :rat-number 11}
-- Failed to map                             -- {:station "cortina", :ltb-harting 0, :paddle-number 114, :ltb-num+channel {:board 11, :ch 8}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 14, :paddle-end :A, :rb-harting 0, :rat-number 11}
-- Failed to map                             -- {:station "cortina", :ltb-harting 0, :paddle-number 115, :ltb-num+channel {:board 11, :ch 6}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 14, :paddle-end :A, :rb-harting 0, :rat-number 11}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 116, :ltb-num+channel {:board 7, :ch 2}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 14, :paddle-end :A, :rb-harting 1, :rat-number 7}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 117, :ltb-num+channel {:board 7, :ch 4}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 14, :paddle-end :A, :rb-harting 1, :rat-number 7}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 118, :ltb-num+channel {:board 7, :ch 6}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 14, :paddle-end :A, :rb-harting 1, :rat-number 7}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 119, :ltb-num+channel {:board 20, :ch 16}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 15, :paddle-end :A, :rb-harting 4, :rat-number 20}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 120, :ltb-num+channel {:board 20, :ch 14}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 15, :paddle-end :A, :rb-harting 4, :rat-number 20}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 121, :ltb-num+channel {:board 20, :ch 12}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 15, :paddle-end :A, :rb-harting 4, :rat-number 20}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 122, :ltb-num+channel {:board 20, :ch 10}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 15, :paddle-end :A, :rb-harting 4, :rat-number 20}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 123, :ltb-num+channel {:board 20, :ch 8}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 15, :paddle-end :A, :rb-harting 4, :rat-number 20}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 124, :ltb-num+channel {:board 20, :ch 6}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 15, :paddle-end :A, :rb-harting 4, :rat-number 20}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 125, :ltb-num+channel {:board 20, :ch 4}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 15, :paddle-end :A, :rb-harting 4, :rat-number 20}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 126, :ltb-num+channel {:board 20, :ch 2}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 15, :paddle-end :A, :rb-harting 4, :rat-number 20}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 127, :ltb-num+channel {:board 13, :ch 16}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 15, :paddle-end :A, :rb-harting 2, :rat-number 13}
-- Failed to map                             -- {:station "cortina", :ltb-harting 0, :paddle-number 128, :ltb-num+channel {:board 11, :ch 2}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 15, :paddle-end :A, :rb-harting 0, :rat-number 11}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 129, :ltb-num+channel {:board 15, :ch 2}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 16, :paddle-end :A, :rb-harting 4, :rat-number 15}
-- Failed to map                             -- {:station "cortina", :ltb-harting 4, :paddle-number 130, :ltb-num+channel {:board 15, :ch 4}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 16, :paddle-end :A, :rb-harting 4, :rat-number 15}
-- Failed to map                             -- {:station "cortina", :ltb-harting 3, :paddle-number 131, :ltb-num+channel {:board 14, :ch 2}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 16, :paddle-end :A, :rb-harting 3, :rat-number 14}
-- Failed to map                             -- {:station "cortina", :ltb-harting 3, :paddle-number 132, :ltb-num+channel {:board 14, :ch 4}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 16, :paddle-end :A, :rb-harting 3, :rat-number 14}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 133, :ltb-num+channel {:board 13, :ch 8}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 16, :paddle-end :A, :rb-harting 2, :rat-number 13}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 134, :ltb-num+channel {:board 13, :ch 10}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 16, :paddle-end :A, :rb-harting 2, :rat-number 13}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 135, :ltb-num+channel {:board 13, :ch 12}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 16, :paddle-end :A, :rb-harting 2, :rat-number 13}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 136, :ltb-num+channel {:board 17, :ch 16}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 16, :paddle-end :A, :rb-harting 1, :rat-number 17}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 137, :ltb-num+channel {:board 17, :ch 14}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 16, :paddle-end :A, :rb-harting 1, :rat-number 17}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 138, :ltb-num+channel {:board 17, :ch 12}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 16, :paddle-end :A, :rb-harting 1, :rat-number 17}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 139, :ltb-num+channel {:board 18, :ch 2}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 17, :paddle-end :A, :rb-harting 2, :rat-number 18}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 140, :ltb-num+channel {:board 18, :ch 4}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 17, :paddle-end :A, :rb-harting 2, :rat-number 18}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 141, :ltb-num+channel {:board 18, :ch 6}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 17, :paddle-end :A, :rb-harting 2, :rat-number 18}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 142, :ltb-num+channel {:board 18, :ch 8}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 17, :paddle-end :A, :rb-harting 2, :rat-number 18}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 143, :ltb-num+channel {:board 18, :ch 10}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 17, :paddle-end :A, :rb-harting 2, :rat-number 18}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 144, :ltb-num+channel {:board 18, :ch 12}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 17, :paddle-end :A, :rb-harting 2, :rat-number 18}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 145, :ltb-num+channel {:board 18, :ch 14}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 17, :paddle-end :A, :rb-harting 2, :rat-number 18}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 146, :ltb-num+channel {:board 18, :ch 16}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 17, :paddle-end :A, :rb-harting 2, :rat-number 18}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 147, :ltb-num+channel {:board 17, :ch 2}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 17, :paddle-end :A, :rb-harting 1, :rat-number 17}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 148, :ltb-num+channel {:board 7, :ch 16}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 17, :paddle-end :A, :rb-harting 1, :rat-number 7}
-- Failed to map                             -- {:station "cortina", :ltb-harting 0, :paddle-number 149, :ltb-num+channel {:board 11, :ch 12}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 18, :paddle-end :A, :rb-harting 0, :rat-number 11}
-- Failed to map                             -- {:station "cortina", :ltb-harting 0, :paddle-number 150, :ltb-num+channel {:board 11, :ch 14}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 18, :paddle-end :A, :rb-harting 0, :rat-number 11}
-- Failed to map                             -- {:station "cortina", :ltb-harting 0, :paddle-number 151, :ltb-num+channel {:board 11, :ch 16}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 18, :paddle-end :A, :rb-harting 0, :rat-number 11}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 152, :ltb-num+channel {:board 13, :ch 1}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 19, :paddle-end :A, :rb-harting 2, :rat-number 13}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 153, :ltb-num+channel {:board 13, :ch 3}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 19, :paddle-end :A, :rb-harting 2, :rat-number 13}
-- Failed to map                             -- {:station "cortina", :ltb-harting 2, :paddle-number 154, :ltb-num+channel {:board 13, :ch 5}, :rb-num+channel :N/A, :dsi-slot 3, :panel-number 19, :paddle-end :A, :rb-harting 2, :rat-number 13}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 155, :ltb-num+channel {:board 17, :ch 5}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 20, :paddle-end :A, :rb-harting 1, :rat-number 17}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 156, :ltb-num+channel {:board 17, :ch 7}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 20, :paddle-end :A, :rb-harting 1, :rat-number 17}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 157, :ltb-num+channel {:board 17, :ch 9}, :rb-num+channel :N/A, :dsi-slot 4, :panel-number 20, :paddle-end :A, :rb-harting 1, :rat-number 17}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 158, :ltb-num+channel {:board 7, :ch 8}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 21, :paddle-end :A, :rb-harting 1, :rat-number 7}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 159, :ltb-num+channel {:board 7, :ch 10}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 21, :paddle-end :A, :rb-harting 1, :rat-number 7}
-- Failed to map                             -- {:station "cortina", :ltb-harting 1, :paddle-number 160, :ltb-num+channel {:board 7, :ch 12}, :rb-num+channel :N/A, :dsi-slot 2, :panel-number 21, :paddle-end :A, :rb-harting 1, :rat-number 7}
  --END: autoinsert mapping

end behavioral;
