`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/29/2022 11:09:42 AM
// Design Name: 
// Module Name: trenzLTproto
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`define PULSE_STEP 1

module
trenzLTproto
   #(parameter GLOBAL_DATE = 0,
     parameter GLOBAL_TIME = 0,
     parameter GLOBAL_VER  = 0,
     parameter GLOBAL_SHA  = 0
     )(
    input       CLK1,

    input [2:0] DISC_A,
    input [2:0] DISC_B,
    input [2:0] DISC_C,
    input [2:0] DISC_D,
    
    input [2:0] DISC_E,
    input [2:0] DISC_F,
    input [2:0] DISC_G,
    input [2:0] DISC_H,
    
    input [2:0] DISC_I,
    input [2:0] DISC_J,
    input [2:0] DISC_K,
    input [2:0] DISC_L,
    
    input [2:0] DISC_M,
    input [2:0] DISC_N,
    input [2:0] DISC_O,
    input [2:0] DISC_P,

    inout       scl, // trenz pin 10 j1, B35_L13_P, F4
    inout       sda, // trenz pin 12 j1, B35_L12_P, E3

    output      LEDgreen,
    
    output      TRIG_OUT_0,
    output      TRIG_OUT_1
    );
    
        
    wire [2:0] thrA;
    wire [2:0] thrB;
    wire [2:0] thrC;
    wire [2:0] thrD;
    
    wire [2:0] thrE;
    wire [2:0] thrF;
    wire [2:0] thrG;
    wire [2:0] thrH;
    
    wire [2:0] thrI;
    wire [2:0] thrJ;
    wire [2:0] thrK;
    wire [2:0] thrL;
    
    wire [2:0] thrM;
    wire [2:0] thrN;
    wire [2:0] thrO;
    wire [2:0] thrP;
    
    
    wire [1:0] bitoutA;
    wire [1:0] bitoutB;
    wire [1:0] bitoutC;
    wire [1:0] bitoutD;
    
    wire [1:0] bitoutE;
    wire [1:0] bitoutF;
    wire [1:0] bitoutG;
    wire [1:0] bitoutH;
    
    
    
    
    reg trigRaw;
    wire tirgDel;
    
    //******swap the 9 and 13 bit version as needed depending on the output format 
    reg [8:0] dataLow;
    //reg [12:0] dataLow;
    reg [8:0] dataHigh;
    //reg [12:0] dataHigh;
    
    
    //turn on the green LED
    assign LEDgreen = 1'b1;   
    
    
    //these are for testing (be sure to disable the regular TRIG_OUT assignments
    //assign TRIG_OUT_0 = DISC_H[0];
    //assign TRIG_OUT_1 = trigDel;
    
    
    //200MHz clock automatically generated by the IP clock wizard
    //CLK2 is the 200MHz clock
    //second argument is 'reset' for the clock, just set to 0 to disable
    //locked is true if the clocks phases are locked
    //final argument is the system (100MHz) clock as input (CLK1)
    clk_wiz_0 ck (CLK2, 0, locked, CLK1);
    
    //these lines set up the individual triggers for each channel and threshold
    //the 200MHz CLK2 is used, so each clock cycle is 5ns
    //******************CLOCK CYCLES START AT 1*******************************
    //.fallingEdge is the where the falling edge is (in clock cycles)
    //.dt is the 'dead time' where the channel/threshold can not trigger again (in clock cycles)
    setreg rA0 (.clk(CLK2), .sig(DISC_A[0]), .fallingEdge(20), .dt(60), .line(thrA[0]));
    setreg rA1 (.clk(CLK2), .sig(DISC_A[1]), .fallingEdge(20), .dt(60), .line(thrA[1]));
    setreg rA2 (.clk(CLK2), .sig(DISC_A[2]), .fallingEdge(20), .dt(60), .line(thrA[2]));
    
    setreg rB0 (.clk(CLK2), .sig(DISC_B[0]), .fallingEdge(20), .dt(60), .line(thrB[0]));
    setreg rB1 (.clk(CLK2), .sig(DISC_B[1]), .fallingEdge(20), .dt(60), .line(thrB[1]));
    setreg rB2 (.clk(CLK2), .sig(DISC_B[2]), .fallingEdge(20), .dt(60), .line(thrB[2]));
    
    setreg rC0 (.clk(CLK2), .sig(DISC_C[0]), .fallingEdge(20), .dt(60), .line(thrC[0]));
    setreg rC1 (.clk(CLK2), .sig(DISC_C[1]), .fallingEdge(20), .dt(60), .line(thrC[1]));
    setreg rC2 (.clk(CLK2), .sig(DISC_C[2]), .fallingEdge(20), .dt(60), .line(thrC[2]));
    
    setreg rD0 (.clk(CLK2), .sig(DISC_D[0]), .fallingEdge(20), .dt(60), .line(thrD[0]));
    setreg rD1 (.clk(CLK2), .sig(DISC_D[1]), .fallingEdge(20), .dt(60), .line(thrD[1]));
    setreg rD2 (.clk(CLK2), .sig(DISC_D[2]), .fallingEdge(20), .dt(60), .line(thrD[2]));
    
    
    setreg rE0 (.clk(CLK2), .sig(DISC_E[0]), .fallingEdge(20), .dt(60), .line(thrE[0]));
    setreg rE1 (.clk(CLK2), .sig(DISC_E[1]), .fallingEdge(20), .dt(60), .line(thrE[1]));
    setreg rE2 (.clk(CLK2), .sig(DISC_E[2]), .fallingEdge(20), .dt(60), .line(thrE[2]));
    
    setreg rF0 (.clk(CLK2), .sig(DISC_F[0]), .fallingEdge(20), .dt(60), .line(thrF[0]));
    setreg rF1 (.clk(CLK2), .sig(DISC_F[1]), .fallingEdge(20), .dt(60), .line(thrF[1]));
    setreg rF2 (.clk(CLK2), .sig(DISC_F[2]), .fallingEdge(20), .dt(60), .line(thrF[2]));
    
    setreg rG0 (.clk(CLK2), .sig(DISC_G[0]), .fallingEdge(20), .dt(60), .line(thrG[0]));
    setreg rG1 (.clk(CLK2), .sig(DISC_G[1]), .fallingEdge(20), .dt(60), .line(thrG[1]));
    setreg rG2 (.clk(CLK2), .sig(DISC_G[2]), .fallingEdge(20), .dt(60), .line(thrG[2]));
    
    //setregClocked rH0 (.clk(CLK2), .sig(DISC_H[0]), .fallingEdge(20), .dt(60), .line(thrH[0]));
    //setregClocked rH1 (.clk(CLK2), .sig(DISC_H[1]), .fallingEdge(20), .dt(60), .line(thrH[1]));
    //setregClocked rH2 (.clk(CLK2), .sig(DISC_H[2]), .fallingEdge(20), .dt(60), .line(thrH[2]));
    
    setreg rH0 (.clk(CLK2), .sig(DISC_H[0]), .fallingEdge(20), .dt(60), .line(thrH[0]));
    setreg rH1 (.clk(CLK2), .sig(DISC_H[1]), .fallingEdge(20), .dt(60), .line(thrH[1]));
    setreg rH2 (.clk(CLK2), .sig(DISC_H[2]), .fallingEdge(20), .dt(60), .line(thrH[2]));
    
    
    setreg rI0 (.clk(CLK2), .sig(DISC_I[0]), .fallingEdge(20), .dt(60), .line(thrI[0]));
    setreg rI1 (.clk(CLK2), .sig(DISC_I[1]), .fallingEdge(20), .dt(60), .line(thrI[1]));
    setreg rI2 (.clk(CLK2), .sig(DISC_I[2]), .fallingEdge(20), .dt(60), .line(thrI[2]));
    
    setreg rJ0 (.clk(CLK2), .sig(DISC_J[0]), .fallingEdge(20), .dt(60), .line(thrJ[0]));
    setreg rJ1 (.clk(CLK2), .sig(DISC_J[1]), .fallingEdge(20), .dt(60), .line(thrJ[1]));
    setreg rJ2 (.clk(CLK2), .sig(DISC_J[2]), .fallingEdge(20), .dt(60), .line(thrJ[2]));
    
    setreg rK0 (.clk(CLK2), .sig(DISC_K[0]), .fallingEdge(20), .dt(60), .line(thrK[0]));
    setreg rK1 (.clk(CLK2), .sig(DISC_K[1]), .fallingEdge(20), .dt(60), .line(thrK[1]));
    setreg rK2 (.clk(CLK2), .sig(DISC_K[2]), .fallingEdge(20), .dt(60), .line(thrK[2]));
    
    setreg rL0 (.clk(CLK2), .sig(DISC_L[0]), .fallingEdge(20), .dt(60), .line(thrL[0]));
    setreg rL1 (.clk(CLK2), .sig(DISC_L[1]), .fallingEdge(20), .dt(60), .line(thrL[1]));
    setreg rL2 (.clk(CLK2), .sig(DISC_L[2]), .fallingEdge(20), .dt(60), .line(thrL[2]));
    
    
    setreg rM0 (.clk(CLK2), .sig(DISC_M[0]), .fallingEdge(20), .dt(60), .line(thrM[0]));
    setreg rM1 (.clk(CLK2), .sig(DISC_M[1]), .fallingEdge(20), .dt(60), .line(thrM[1]));
    setreg rM2 (.clk(CLK2), .sig(DISC_M[2]), .fallingEdge(20), .dt(60), .line(thrM[2]));
    
    setreg rN0 (.clk(CLK2), .sig(DISC_N[0]), .fallingEdge(20), .dt(60), .line(thrN[0]));
    setreg rN1 (.clk(CLK2), .sig(DISC_N[1]), .fallingEdge(20), .dt(60), .line(thrN[1]));
    setreg rN2 (.clk(CLK2), .sig(DISC_N[2]), .fallingEdge(20), .dt(60), .line(thrN[2]));
    
    setreg rO0 (.clk(CLK2), .sig(DISC_O[0]), .fallingEdge(20), .dt(60), .line(thrO[0]));
    setreg rO1 (.clk(CLK2), .sig(DISC_O[1]), .fallingEdge(20), .dt(60), .line(thrO[1]));
    setreg rO2 (.clk(CLK2), .sig(DISC_O[2]), .fallingEdge(20), .dt(60), .line(thrO[2]));
    
    setreg rP0 (.clk(CLK2), .sig(DISC_P[0]), .fallingEdge(20), .dt(60), .line(thrP[0]));
    setreg rP1 (.clk(CLK2), .sig(DISC_P[1]), .fallingEdge(20), .dt(60), .line(thrP[1]));
    setreg rP2 (.clk(CLK2), .sig(DISC_P[2]), .fallingEdge(20), .dt(60), .line(thrP[2]));
    
    //set a delay and pulse width on the trigger (formed below from thr0's)
    //data starts getting sent after the falling edge of the trigger
    //delay falling edge of trig signal enough to capture thr2 at high amplitude
    //some delay on falling edge seems necessary to ensure higher thresholds are captured correctly
    setregClocked tr (.clk(CLK2), .sig(trigRaw), .fallingEdge(5), .dt(15), .line(trigDel));
    
    
    
    //these will set the bit combinations if we are using the 9-bit output version 
    makeBitNC bA (.thr0(thrA[0] | thrB[0]), .thr1(thrA[1] | thrB[1]), .thr2(thrA[2] | thrB[2]), .bitout(bitoutA));
    makeBitNC bB (.thr0(thrC[0] | thrD[0]), .thr1(thrC[1] | thrD[1]), .thr2(thrC[2] | thrD[2]), .bitout(bitoutB));
    makeBitNC bC (.thr0(thrE[0] | thrF[0]), .thr1(thrE[1] | thrF[1]), .thr2(thrE[2] | thrF[2]), .bitout(bitoutC));
    makeBitNC bD (.thr0(thrG[0] | thrH[0]), .thr1(thrG[1] | thrH[1]), .thr2(thrG[2] | thrH[2]), .bitout(bitoutD));
    
    makeBitNC bE (.thr0(thrI[0] | thrJ[0]), .thr1(thrI[1] | thrJ[1]), .thr2(thrI[2] | thrJ[2]), .bitout(bitoutE));
    makeBitNC bF (.thr0(thrK[0] | thrL[0]), .thr1(thrK[1] | thrL[1]), .thr2(thrK[2] | thrL[2]), .bitout(bitoutF));
    makeBitNC bG (.thr0(thrM[0] | thrN[0]), .thr1(thrM[1] | thrN[1]), .thr2(thrM[2] | thrN[2]), .bitout(bitoutG));
    makeBitNC bH (.thr0(thrO[0] | thrP[0]), .thr1(thrO[1] | thrP[1]), .thr2(thrO[2] | thrP[2]), .bitout(bitoutH));

    
    
    always @ * begin
        //dataLow = {1'b1, thrA[0] | thrI[0], thrB[0] | thrJ[0] ,thrC[0] | thrK[0] ,thrD[0] | thrL[0] ,thrE[0] | thrM[0], thrF[0] | thrN[0],thrG[0] | thrO[0] , thrH[0] | thrP[0]};
        //dataMid = {1'b1, thrA[1] | thrI[1], thrB[1] | thrJ[1] ,thrC[1] | thrK[1] ,thrD[1] | thrL[1] ,thrE[1] | thrM[1], thrF[1] | thrN[1],thrG[1] | thrO[1] , thrH[1] | thrP[1]};
        //dataHigh = {1'b1, thrA[2] | thrI[2], thrB[2] | thrJ[2] ,thrC[2] | thrK[2] ,thrD[2] | thrL[2] ,thrE[2] | thrM[2], thrF[2] | thrN[2],thrG[2] | thrO[2] , thrH[2] | thrP[2]};
        //veto = (thrA[2] | thrB[2] | thrC[2] | thrD[2] | thrE[2] | thrF[2] | thrG[2] | thrH[2] | thrI[2] | thrJ[2] | thrK[2] | thrL[2] | thrM[2] | thrN[2] | thrO[2] | thrP[2]);
        
        //13 bit each link thr2-first version, format is:
        //dataLow = START bit+thr0 bitmask (8 bits)+thr1 bitmmask (first 4)
        //dataHigh = START bit+thr2 bitmaks (8 bits) + thr1 bitmask (last 4 bits)
        //uncomment the following two lines
        //dataLow  = {1'b1, thrA[0] | thrI[0], thrB[0] | thrJ[0] ,thrC[0] | thrK[0] ,thrD[0] | thrL[0] ,thrE[0] | thrM[0], thrF[0] | thrN[0],thrG[0] | thrO[0] , thrH[0] | thrP[0], thrA[1] | thrI[1], thrB[1] | thrJ[1] ,thrC[1] | thrK[1] ,thrD[1] | thrL[1] };
        //dataHigh = {1'b1, thrA[2] | thrI[2], thrB[2] | thrJ[2] ,thrC[2] | thrK[2] ,thrD[2] | thrL[2] ,thrE[2] | thrM[2], thrF[2] | thrN[2],thrG[2] | thrO[2] , thrH[2] | thrP[2], thrE[1] | thrM[1], thrF[1] | thrN[1],thrG[1] | thrO[1] , thrH[1] | thrP[1] };
        
        //13 bit each link thr1-first version, format is:
        //dataLow  = START bit+thr0 bitmask (8 bits) + thr2 bitmmask (first 4)
        //dataHigh = START bit+thr1 bitmask (8 bits) + thr2 bitmask (last 4 bits)
        //uncomment the following two lines
        //dataLow  = {1'b1, thrA[0] | thrI[0], thrB[0] | thrJ[0] ,thrC[0] | thrK[0] ,thrD[0] | thrL[0] ,thrE[0] | thrM[0], thrF[0] | thrN[0],thrG[0] | thrO[0] , thrH[0] | thrP[0], thrA[2] | thrI[2], thrB[2] | thrJ[2], thrC[2] | thrK[2], thrD[2] | thrL[2] };
        //dataHigh = {1'b1, thrA[1] | thrI[1], thrB[1] | thrJ[1] ,thrC[1] | thrK[1] ,thrD[1] | thrL[1] ,thrE[1] | thrM[1], thrF[1] | thrN[1],thrG[1] | thrO[1] , thrH[1] | thrP[1], thrE[2] | thrM[2], thrF[2] | thrN[2], thrG[2] | thrO[2], thrH[2] | thrP[2] };
        
        //9 bit each link, each paddle has a two bits available (LINK0, LINK1), truth table is:
        
        //      | no hit| thr0 | thr1 | thr2 
        //----------------------------------
        // bit0 |    0  |  0   |  1   |  1
        // bit1 |    0  |  1   |  0   |  1
        
        //dataLow  = START bit +paddles bit 0 (9 bits total)
        //dataHigh = START bit +paddles bit 1 (9 bits total)
        //bitOut 
        
        dataLow  = {1'b1, bitoutA[0], bitoutB[0], bitoutC[0], bitoutD[0], bitoutE[0], bitoutF[0], bitoutG[0], bitoutH[0]};
        dataHigh = {1'b1, bitoutA[1], bitoutB[1], bitoutC[1], bitoutD[1], bitoutE[1], bitoutF[1], bitoutG[1], bitoutH[1]};
        
        
        //trigger formation happens here (this will start the trigger sending process)
        trigRaw = (thrA[0] | thrB[0] | thrC[0] | thrD[0] | thrE[0] | thrF[0] | thrG[0] | thrH[0] | thrI[0] | thrJ[0] | thrK[0] | thrL[0] | thrM[0] | thrN[0] | thrO[0] | thrP[0]);

    end
    
    
    //this is for the trigger package types with 9 bits
    shiftPISO9 s0 (.clk(CLK2), .trig(trigDel), .data(dataLow), .line(TRIG_OUT_0) );
    shiftPISO9 s1 (.clk(CLK2), .trig(trigDel), .data(dataHigh), .line(TRIG_OUT_1) );

    //this is for the trigger package types with 13 bits 
    //shiftPISO13 s0 (.clk(CLK2), .trig(trigDel), .data(dataLow), .line(TRIG_OUT_0) );
    //shiftPISO13 s1 (.clk(CLK2), .trig(trigDel), .data(dataHigh), .line(TRIG_OUT_1) );   


   // `define I2C_ADDRESS 7'h3c
   i2cSlave u_i2cSlave
     (
      .clk(CLK2),
      .rst(!locked),
      .sda(sda),
      .scl(scl),
      .myReg0(),
      .myReg1(),
      .myReg2(),
      .myReg3(),
      .myReg4(GLOBAL_SHA[7:0]),
      .myReg5(GLOBAL_SHA[15:8]),
      .myReg6(GLOBAL_SHA[23:16]),
      .myReg7(GLOBAL_SHA[31:24])
      );

endmodule


//taken from PISO shift register example from here https://techmasterplus.com/programs/verilog/verilog-shiftregister.php?i=1
//9 bit version
module shiftPISO9(clk, trig, data, line);
    input clk;
    input trig;
    input [8:0] data;//9 bits, trigger bit plus 8 bits for paddles bitmask
    output reg line;
    
    reg [8:0] tempData;
    reg [3:0] hold_count;
    
     always @ (posedge clk) begin
        if(trig) begin
            tempData<=data;
            end
        else begin
            line<=tempData[8];
            tempData<={tempData[7:0], 1'b0};
            end
        end
endmodule

//taken from PISO shift register example from here https://techmasterplus.com/programs/verilog/verilog-shiftregister.php?i=1
//13 bit version
module shiftPISO13(clk, trig, data, line);
    input clk;
    input trig;
    input [12:0] data;//13 bits, trigger bit plus 12 bits for paddles bitmask
    output reg line;
    
    reg [12:0] tempData;
    reg [3:0] hold_count;
    
     always @ (posedge clk) begin
        if(trig) begin
            tempData<=data;
            end
        else begin
            line<=tempData[12];
            tempData<={tempData[11:0], 1'b0};
            end
        end
endmodule

//this module will set a register high on a non-clocked edge
//clears after a selectable time (in clock cycles)
module setreg(clk, sig, fallingEdge, dt, line);
    input clk;
    input sig;
    input [7:0] fallingEdge;//pulse width in number of clock counts
    input [7:0] dt;//'dead time' where line is blocked from being set to on again
    output reg line;
    
    
    reg clear = 1'b0;
    reg[7:0] count = 8'b0;
    reg hold = 1'b0;
    
    //wire cl;
    //assign cl = clear;
    
    always@ * begin
        line = (sig & !clear) | (hold & !clear);  
        end
    
        
    always@ (posedge clk) begin           
        if(line && count==0) begin //start counting if line is high this clock cycle
            count<=1;
            hold<=1'b1;//this will keep line high until we clear it
            end    
        if(count==fallingEdge) begin//if count reaches the pulse width, set clear high and hold to low
            clear<=1'b1;
            hold<=1'b0;
            end
        if(count==dt) begin //once dt counter is reached, set clear to 0 and reset the counter, so line can be set high again by the next event
            clear<=1'b0;
            count<=0;
            end   
        if(count>0) begin//incirment counter if event has started
            count<=count+1;
            end
        end        
            
endmodule


//this module will set a register high on a clock edge after the input goes high
//user selectable amount of delay to set falling edge and dead time
module setregClocked(clk, sig, fallingEdge, dt, line);
    input clk;
    input sig;
    input [7:0] fallingEdge;//falling edge of output (in clock counts)
    input [7:0] dt;//'dead time' where line is blocked from being set to high again
    output reg line;
    
    
    reg[7:0] count = 8'b0;
    //reg inEvent = 1'b0;
        
    always@ (posedge clk) begin           
        if(sig && count==0) begin //start counting if input signal is high this clock cycle
            count<=1;
            line<=1'b1;//set the output line high
            end
        if(count==fallingEdge) begin//end the pulse ones this count is reached
            line<=1'b0;
            end
        if(count==dt) begin //once 'dead'time counter is reached, reset the counter, new event can now come in
            count<=0;
            end   
        if(count>0) begin//incirment counter if event has started
            count<=count+1;
            end
        end        
            
endmodule

//non-clocked module to set the trigger output bits correctly for a given input
module makeBitNC(thr0, thr1, thr2, bitout);
    input thr0;
    input thr1;
    input thr2;
    output reg [1:0] bitout;
    
    always@ * begin
    
        if(!thr0 && !thr1 && !thr2) begin
            bitout=2'b00;
            end
    
        else if(thr0 && !thr1 && !thr2) begin//threshold 0 only crossed
            bitout=2'b01;
            end
                
        else if(thr1 && !thr2) begin//threshold 1 but not 2 crossed
            bitout=2'b10;
            end
         
        else if(thr2) begin//threshold 2 crossed
            bitout=2'b11;
            end
            
        else begin //something went wrong, this should not happen
            bitout=2'b00;
            end
           
        end//end of always@ * statement 

endmodule




